
module FIR_FILTER2_DW01_add_0 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_1 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_2 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_3 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_4 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_5 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_6 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_7 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_8 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_9 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_10 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_11 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_12 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_13 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_14 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_15 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_30 ( B, SUM, A_31_, A_30_, A_29_, A_28_, A_27_, 
        A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [31:0] B;
  output [31:0] SUM;
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_;

  wire   [31:1] carry;

  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CMPR32X2 U1_2 ( .A(A_2_), .B(B[2]), .C(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_1 ( .A(A_1_), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_29 ( A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, 
        A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, A_3_, A_2_, A_1_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, 
        B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, 
        B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, 
        B_4_, B_3_, B_2_, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, 
        SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_
 );
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_,
         SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_,
         SUM_2_, SUM_1_;

  wire   [31:1] carry;

  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM_31_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFHX2 U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFHX2 U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFHX2 U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFHX2 U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFHX2 U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFHX2 U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFHX2 U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFHX2 U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFHX2 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFHX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFHX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFHX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX2 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_1 ( .A(A_1_), .B(1'b0), .CI(1'b0), .S(SUM_1_) );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(1'b0), .CO(carry[3]), .S(SUM_2_) );
endmodule


module FIR_FILTER2_DW01_add_28 ( A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, 
        A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, A_3_, A_2_, A_1_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, 
        B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, 
        B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, 
        B_4_, B_3_, B_2_, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, 
        SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_
 );
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_,
         SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_,
         SUM_2_, SUM_1_;

  wire   [31:1] carry;

  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM_31_) );
  ADDFXL U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFXL U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  CMPR32X2 U1_8 ( .A(A_8_), .B(B_8_), .C(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  CMPR32X2 U1_7 ( .A(A_7_), .B(B_7_), .C(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFXL U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFHX2 U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFHX4 U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFHX2 U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFHX2 U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFHX4 U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFHX2 U1_1 ( .A(A_1_), .B(1'b0), .CI(1'b0), .S(SUM_1_) );
  ADDFHX2 U1_2 ( .A(A_2_), .B(B_2_), .CI(1'b0), .CO(carry[3]), .S(SUM_2_) );
endmodule


module FIR_FILTER2_DW01_add_27 ( A, SUM, B_31_, B_30_, B_29_, B_28_, B_27_, 
        B_26_, B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, 
        B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_ );
  input [31:0] A;
  output [31:0] SUM;
  input B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;

  wire   [31:1] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B_31_), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_11 ( .A(A[11]), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  CMPR32X2 U1_8 ( .A(A[8]), .B(B_8_), .C(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_24 ( .A(A[24]), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX1 U1_13 ( .A(A[13]), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX1 U1_7 ( .A(A[7]), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_9 ( .A(A[9]), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_10 ( .A(A[10]), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B_1_), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_26 ( A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, 
        A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, A_3_, A_2_, A_1_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, 
        B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, 
        B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, 
        B_4_, B_3_, B_2_, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, 
        SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, 
        SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_
 );
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_,
         SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_,
         SUM_2_, SUM_1_;

  wire   [31:1] carry;

  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM_31_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFHX2 U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFHX2 U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFHX2 U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFHX2 U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFHX2 U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFHX4 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFHX2 U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFHX2 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX2 U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_1 ( .A(A_1_), .B(1'b0), .CI(1'b0), .S(SUM_1_) );
  CMPR32X2 U1_2 ( .A(A_2_), .B(B_2_), .C(1'b0), .CO(carry[3]), .S(SUM_2_) );
endmodule


module FIR_FILTER2_DW01_add_25 ( A, SUM, B_31_, B_30_, B_29_, B_28_, B_27_, 
        B_26_, B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, 
        B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_ );
  input [31:0] A;
  output [31:0] SUM;
  input B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;
  wire   n2, n3, n4, n5;
  wire   [31:1] carry;

  ADDFXL U1_15 ( .A(A[15]), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  XOR3X1 U1_31 ( .A(A[31]), .B(B_31_), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_2 ( .A(A[2]), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_26 ( .A(A[26]), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_6 ( .A(A[6]), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_4 ( .A(A[4]), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_5 ( .A(A[5]), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B_1_), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
  NAND3X1 U3 ( .A(n3), .B(n4), .C(n5), .Y(carry[4]) );
  NAND2X1 U4 ( .A(A[3]), .B(B_3_), .Y(n5) );
  XOR2X1 U5 ( .A(carry[3]), .B(n2), .Y(SUM[3]) );
  XOR2XL U6 ( .A(B_3_), .B(A[3]), .Y(n2) );
  NAND2X2 U7 ( .A(B_3_), .B(carry[3]), .Y(n3) );
  NAND2X2 U8 ( .A(A[3]), .B(carry[3]), .Y(n4) );
endmodule


module FIR_FILTER2_DW01_add_24 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:2] carry;

  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  CMPR32X2 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFHX4 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_23 ( A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, 
        A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, A_3_, A_2_, A_1_, B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, 
        B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, 
        B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, 
        B_4_, B_3_, B_2_, B_1_, SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, 
        SUM_26_, SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, 
        SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, 
        SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, 
        SUM_2_, SUM_1_ );
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_,
         SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_,
         SUM_2_, SUM_1_;

  wire   [31:1] carry;

  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  XOR3X1 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM_31_) );
  ADDFXL U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFXL U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFX1 U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  ADDFX1 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFHX4 U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFHX4 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFHX4 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFHX4 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFX2 U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFXL U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFXL U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFXL U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFHX1 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFX2 U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFX2 U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFHX2 U1_1 ( .A(A_1_), .B(B_1_), .CI(1'b0), .CO(carry[2]), .S(SUM_1_) );
endmodule


module FIR_FILTER2_DW01_add_22 ( B, SUM, A_31_, A_30_, A_29_, A_28_, A_27_, 
        A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [31:0] B;
  output [31:0] SUM;
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_;

  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A_31_), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_8 ( .A(A_8_), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  CMPR32X2 U1_9 ( .A(A_9_), .B(B[9]), .C(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX2 U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_28 ( .A(A_28_), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_25 ( .A(A_25_), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX2 U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  CMPR32X2 U1_18 ( .A(A_18_), .B(B[18]), .C(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX2 U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_1 ( .A(A_1_), .B(B[1]), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_21 ( A, SUM, B_31_, B_30_, B_29_, B_28_, B_27_, 
        B_26_, B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, 
        B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_ );
  input [31:0] A;
  output [31:0] SUM;
  input B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;

  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B_31_), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX1 U1_14 ( .A(A[14]), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX1 U1_15 ( .A(A[15]), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_17 ( .A(A[17]), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  CMPR32X2 U1_27 ( .A(A[27]), .B(B_27_), .C(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX1 U1_13 ( .A(A[13]), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_30 ( .A(A[30]), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B_1_), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_20 ( A, SUM, B_31_, B_30_, B_29_, B_28_, B_27_, 
        B_26_, B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, 
        B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_ );
  input [31:0] A;
  output [31:0] SUM;
  input B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_;

  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A[31]), .B(B_31_), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX1 U1_15 ( .A(A[15]), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_24 ( .A(A[24]), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX1 U1_26 ( .A(A[26]), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  CMPR32X2 U1_2 ( .A(A[2]), .B(B_2_), .C(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CMPR32X2 U1_29 ( .A(A[29]), .B(B_29_), .C(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX2 U1_12 ( .A(A[12]), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  CMPR32X2 U1_27 ( .A(A[27]), .B(B_27_), .C(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX1 U1_21 ( .A(A[21]), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX1 U1_25 ( .A(A[25]), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX1 U1_1 ( .A(A[1]), .B(B_1_), .CI(1'b0), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(1'b0), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_19 ( B, SUM, A_31_, A_30_, A_29_, A_28_, A_27_, 
        A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, A_3_, A_2_, A_1_ );
  input [31:0] B;
  output [31:0] SUM;
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [31:2] carry;

  XOR3X1 U1_31 ( .A(A_31_), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_22 ( .A(A_22_), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_3 ( .A(A_3_), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFHX4 U1_29 ( .A(A_29_), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_27 ( .A(A_27_), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_4 ( .A(A_4_), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFHX4 U1_13 ( .A(A_13_), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX4 U1_7 ( .A(A_7_), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A_6_), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A_5_), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX2 U1_11 ( .A(A_11_), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  CMPR32X2 U1_2 ( .A(A_2_), .B(B[2]), .C(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFHX4 U1_30 ( .A(A_30_), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_26 ( .A(A_26_), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_24 ( .A(A_24_), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  CMPR32X2 U1_25 ( .A(A_25_), .B(B[25]), .C(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_23 ( .A(A_23_), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  CLKINVX6 U1 ( .A(n10), .Y(carry[2]) );
  XOR2X4 U2 ( .A(B[1]), .B(A_1_), .Y(SUM[1]) );
  XOR2X1 U3 ( .A(B[0]), .B(1'b0), .Y(SUM[0]) );
  XOR2X4 U5 ( .A(B[28]), .B(A_28_), .Y(n11) );
  XOR2XL U6 ( .A(carry[12]), .B(n6), .Y(SUM[12]) );
  XOR2XL U7 ( .A(A_12_), .B(B[12]), .Y(n6) );
  NAND3X1 U8 ( .A(n3), .B(n4), .C(n5), .Y(carry[9]) );
  XOR2X1 U9 ( .A(carry[8]), .B(n2), .Y(SUM[8]) );
  XOR2X1 U10 ( .A(A_8_), .B(B[8]), .Y(n2) );
  NAND2X1 U11 ( .A(B[12]), .B(carry[12]), .Y(n8) );
  NAND2X1 U12 ( .A(A_28_), .B(carry[28]), .Y(n13) );
  XOR2X1 U13 ( .A(carry[28]), .B(n11), .Y(SUM[28]) );
  NAND2X1 U14 ( .A(A_8_), .B(carry[8]), .Y(n3) );
  NAND2X1 U15 ( .A(B[8]), .B(carry[8]), .Y(n4) );
  NAND2X1 U16 ( .A(B[8]), .B(A_8_), .Y(n5) );
  NAND2X2 U17 ( .A(A_12_), .B(carry[12]), .Y(n7) );
  NAND2X4 U18 ( .A(B[12]), .B(A_12_), .Y(n9) );
  NAND3X6 U19 ( .A(n7), .B(n8), .C(n9), .Y(carry[13]) );
  NAND2X1 U20 ( .A(A_1_), .B(B[1]), .Y(n10) );
  NAND2X4 U21 ( .A(B[28]), .B(carry[28]), .Y(n12) );
  NAND2X4 U22 ( .A(A_28_), .B(B[28]), .Y(n14) );
  NAND3X4 U23 ( .A(n12), .B(n13), .C(n14), .Y(carry[29]) );
endmodule


module FIR_FILTER2_DW01_add_18 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1;
  wire   [31:2] carry;

  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  CMPR32X2 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  CMPR32X2 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFHX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_17 ( A, B, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [31:2] carry;

  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  CMPR32X2 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  CMPR32X2 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFHX4 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX4 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFHX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX4 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX4 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  XOR3X1 U1 ( .A(A[2]), .B(B[2]), .C(carry[2]), .Y(SUM[2]) );
  XOR3X1 U2 ( .A(B[6]), .B(carry[6]), .C(A[6]), .Y(SUM[6]) );
  AND2X2 U3 ( .A(B[0]), .B(A[0]), .Y(n1) );
  NAND2XL U4 ( .A(A[6]), .B(B[6]), .Y(n2) );
  NAND2XL U5 ( .A(carry[6]), .B(B[6]), .Y(n3) );
  NAND2XL U6 ( .A(carry[6]), .B(A[6]), .Y(n4) );
  NAND3X1 U7 ( .A(n2), .B(n3), .C(n4), .Y(carry[7]) );
  XOR3X2 U8 ( .A(B[4]), .B(carry[4]), .C(A[4]), .Y(SUM[4]) );
  NAND2XL U9 ( .A(A[4]), .B(B[4]), .Y(n5) );
  NAND2XL U10 ( .A(carry[4]), .B(B[4]), .Y(n6) );
  NAND2XL U11 ( .A(carry[4]), .B(A[4]), .Y(n7) );
  NAND3X1 U12 ( .A(n5), .B(n6), .C(n7), .Y(carry[5]) );
  NAND2XL U13 ( .A(carry[2]), .B(A[2]), .Y(n8) );
  NAND2XL U14 ( .A(B[2]), .B(A[2]), .Y(n9) );
  NAND2XL U15 ( .A(B[2]), .B(carry[2]), .Y(n10) );
  NAND3X1 U16 ( .A(n8), .B(n9), .C(n10), .Y(carry[3]) );
  XOR2X1 U17 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW01_add_16 ( A, B, SUM_31_, SUM_30_, SUM_29_, SUM_28_, 
        SUM_27_, SUM_26_, SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, 
        SUM_19_, SUM_18_, SUM_17_, SUM_16_ );
  input [31:0] A;
  input [31:0] B;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [31:16] carry;

  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM_29_) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM_26_) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM_31_) );
  ADDFX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM_25_) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM_27_) );
  CMPR32X2 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM_28_) );
  ADDFX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM_23_) );
  ADDFX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM_22_) );
  ADDFX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  ADDFX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM_30_) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM_24_) );
  OAI2BB1X2 U1 ( .A0N(n6), .A1N(A[13]), .B0(n7), .Y(n4) );
  OAI21X1 U2 ( .A0(A[6]), .A1(n20), .B0(B[6]), .Y(n21) );
  OAI21X4 U3 ( .A0(A[14]), .A1(n4), .B0(B[14]), .Y(n5) );
  OAI2BB1X4 U4 ( .A0N(n4), .A1N(A[14]), .B0(n5), .Y(n3) );
  OAI21X1 U5 ( .A0(A[4]), .A1(n24), .B0(B[4]), .Y(n25) );
  BUFX4 U6 ( .A(A[15]), .Y(n1) );
  OAI2BB1X4 U7 ( .A0N(n22), .A1N(A[5]), .B0(n23), .Y(n20) );
  OAI21X4 U8 ( .A0(A[5]), .A1(n22), .B0(B[5]), .Y(n23) );
  OAI2BB1X4 U9 ( .A0N(n18), .A1N(A[7]), .B0(n19), .Y(n16) );
  OAI21X4 U10 ( .A0(A[7]), .A1(n18), .B0(B[7]), .Y(n19) );
  OAI21X2 U11 ( .A0(A[3]), .A1(n26), .B0(B[3]), .Y(n27) );
  OAI2BB1X2 U12 ( .A0N(n28), .A1N(A[2]), .B0(n29), .Y(n26) );
  OAI2BB1X4 U13 ( .A0N(n26), .A1N(A[3]), .B0(n27), .Y(n24) );
  OAI2BB1X1 U14 ( .A0N(n20), .A1N(A[6]), .B0(n21), .Y(n18) );
  OAI2BB1X1 U15 ( .A0N(n14), .A1N(A[9]), .B0(n15), .Y(n12) );
  OAI21X1 U16 ( .A0(A[9]), .A1(n14), .B0(B[9]), .Y(n15) );
  OAI2BB1X1 U17 ( .A0N(n16), .A1N(A[8]), .B0(n17), .Y(n14) );
  OAI21X1 U18 ( .A0(A[8]), .A1(n16), .B0(B[8]), .Y(n17) );
  OAI2BB1X2 U19 ( .A0N(n8), .A1N(A[12]), .B0(n9), .Y(n6) );
  OAI21X1 U20 ( .A0(A[11]), .A1(n10), .B0(B[11]), .Y(n11) );
  OAI2BB1X1 U21 ( .A0N(n12), .A1N(A[10]), .B0(n13), .Y(n10) );
  OAI21X2 U22 ( .A0(A[10]), .A1(n12), .B0(B[10]), .Y(n13) );
  OAI21X4 U23 ( .A0(A[13]), .A1(n6), .B0(B[13]), .Y(n7) );
  OAI21X4 U24 ( .A0(A[12]), .A1(n8), .B0(B[12]), .Y(n9) );
  OAI2BB1X1 U25 ( .A0N(n24), .A1N(A[4]), .B0(n25), .Y(n22) );
  OAI21X1 U26 ( .A0(A[2]), .A1(n28), .B0(B[2]), .Y(n29) );
  AO21X4 U27 ( .A0(n3), .A1(n1), .B0(n2), .Y(carry[16]) );
  OA21X4 U28 ( .A0(n1), .A1(n3), .B0(B[15]), .Y(n2) );
  OAI2BB1X1 U29 ( .A0N(A[1]), .A1N(B[1]), .B0(n30), .Y(n28) );
  OAI211X1 U30 ( .A0(A[1]), .A1(B[1]), .B0(A[0]), .C0(B[0]), .Y(n30) );
  OAI2BB1X1 U31 ( .A0N(n10), .A1N(A[11]), .B0(n11), .Y(n8) );
endmodule


module FIR_FILTER2_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module FIR_FILTER2_DW_mult_uns_15 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n157, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182;

  ADDFXL U16 ( .A(a_15_), .B(n168), .CI(n12), .CO(n11), .S(product_22_) );
  ADDFXL U17 ( .A(n33), .B(a_14_), .CI(n13), .CO(n12), .S(product_21_) );
  ADDFXL U18 ( .A(n34), .B(n35), .CI(n14), .CO(n13), .S(product_20_) );
  ADDFXL U19 ( .A(n37), .B(n36), .CI(n15), .CO(n14), .S(product_19_) );
  ADDFXL U20 ( .A(n39), .B(n38), .CI(n16), .CO(n15), .S(product_18_) );
  ADDFXL U21 ( .A(n41), .B(n40), .CI(n17), .CO(n16), .S(product_17_) );
  ADDFXL U22 ( .A(n43), .B(n42), .CI(n18), .CO(n17), .S(product_16_) );
  ADDFXL U23 ( .A(n44), .B(n45), .CI(n19), .CO(n18), .S(product_15_) );
  ADDFXL U24 ( .A(n46), .B(n47), .CI(n20), .CO(n19), .S(product_14_) );
  ADDFXL U25 ( .A(n48), .B(n49), .CI(n21), .CO(n20), .S(product_13_) );
  ADDFXL U26 ( .A(n50), .B(n51), .CI(n22), .CO(n21), .S(product_12_) );
  ADDFXL U27 ( .A(n52), .B(n53), .CI(n23), .CO(n22), .S(product_11_) );
  ADDFXL U28 ( .A(n54), .B(n55), .CI(n24), .CO(n23), .S(product_10_) );
  ADDFXL U29 ( .A(n56), .B(n57), .CI(n25), .CO(n24), .S(product_9_) );
  ADDFXL U30 ( .A(n58), .B(n59), .CI(n26), .CO(n25), .S(product_8_) );
  ADDFXL U31 ( .A(n60), .B(a_2_), .CI(n27), .CO(n26), .S(product_7_) );
  ADDFXL U32 ( .A(a_1_), .B(n177), .CI(n28), .CO(n27), .S(product_6_) );
  ADDFXL U33 ( .A(a_0_), .B(n178), .CI(n29), .CO(n28), .S(product_5_) );
  ADDHXL U34 ( .A(n179), .B(n30), .CO(n29), .S(product_4_) );
  ADDHXL U35 ( .A(n180), .B(n31), .CO(n30), .S(product_3_) );
  ADDHXL U36 ( .A(n181), .B(n182), .CO(n31), .S(product_2_) );
  ADDFXL U38 ( .A(n170), .B(n167), .CI(n169), .CO(n33), .S(n34) );
  ADDFXL U39 ( .A(n171), .B(a_12_), .CI(a_14_), .CO(n35), .S(n36) );
  ADDFXL U40 ( .A(n172), .B(a_11_), .CI(a_13_), .CO(n37), .S(n38) );
  ADDFXL U41 ( .A(n173), .B(a_10_), .CI(a_12_), .CO(n39), .S(n40) );
  ADDFXL U42 ( .A(a_15_), .B(a_9_), .CI(a_11_), .CO(n41), .S(n42) );
  ADDFXL U43 ( .A(n174), .B(n168), .CI(a_10_), .CO(n43), .S(n44) );
  ADDFXL U44 ( .A(n175), .B(n169), .CI(a_9_), .CO(n45), .S(n46) );
  ADDFXL U45 ( .A(n176), .B(n170), .CI(a_8_), .CO(n47), .S(n48) );
  ADDFXL U46 ( .A(n177), .B(n171), .CI(a_7_), .CO(n49), .S(n50) );
  ADDFXL U47 ( .A(n178), .B(n172), .CI(a_6_), .CO(n51), .S(n52) );
  ADDFXL U48 ( .A(n179), .B(n173), .CI(a_5_), .CO(n53), .S(n54) );
  ADDFXL U49 ( .A(n180), .B(n174), .CI(a_4_), .CO(n55), .S(n56) );
  ADDFXL U50 ( .A(n181), .B(n175), .CI(a_3_), .CO(n57), .S(n58) );
  INVX3 U73 ( .A(product_28_), .Y(n157) );
  CLKINVX1 U74 ( .A(n11), .Y(product_28_) );
  CLKINVX1 U75 ( .A(n157), .Y(product_23_) );
  CLKINVX1 U76 ( .A(n157), .Y(product_24_) );
  CLKINVX1 U77 ( .A(n157), .Y(product_25_) );
  CLKINVX1 U78 ( .A(n157), .Y(product_26_) );
  CLKINVX1 U79 ( .A(n157), .Y(product_27_) );
  CLKINVX1 U80 ( .A(n157), .Y(product_29_) );
  CLKINVX1 U81 ( .A(n157), .Y(product_30_) );
  CLKINVX1 U82 ( .A(n157), .Y(product_31_) );
  CLKINVX1 U83 ( .A(a_0_), .Y(n182) );
  CLKINVX1 U84 ( .A(a_3_), .Y(n179) );
  CLKINVX1 U85 ( .A(a_4_), .Y(n178) );
  CLKINVX1 U86 ( .A(a_5_), .Y(n177) );
  CLKINVX1 U87 ( .A(a_7_), .Y(n175) );
  CLKINVX1 U88 ( .A(a_2_), .Y(n180) );
  CLKINVX1 U89 ( .A(a_1_), .Y(n181) );
  CLKINVX1 U90 ( .A(a_6_), .Y(n176) );
  CLKINVX1 U91 ( .A(a_9_), .Y(n173) );
  CLKINVX1 U92 ( .A(a_10_), .Y(n172) );
  CLKINVX1 U93 ( .A(a_8_), .Y(n174) );
  CLKINVX1 U94 ( .A(a_11_), .Y(n171) );
  CLKINVX1 U95 ( .A(a_12_), .Y(n170) );
  CLKINVX1 U96 ( .A(a_13_), .Y(n169) );
  CLKINVX1 U97 ( .A(a_14_), .Y(n168) );
  CLKINVX1 U98 ( .A(a_15_), .Y(n167) );
  CLKBUFX3 U99 ( .A(a_0_), .Y(product_1_) );
  XOR2X1 U100 ( .A(n176), .B(a_0_), .Y(n60) );
  NAND2X1 U101 ( .A(a_0_), .B(a_6_), .Y(n59) );
endmodule


module FIR_FILTER2_DW_mult_uns_14 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n148,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172;

  ADDFXL U16 ( .A(a_15_), .B(n159), .CI(n12), .CO(n11), .S(product_22_) );
  ADDFXL U17 ( .A(n160), .B(a_14_), .CI(n13), .CO(n12), .S(product_21_) );
  ADDFXL U18 ( .A(n161), .B(a_13_), .CI(n14), .CO(n13), .S(product_20_) );
  ADDFXL U19 ( .A(n162), .B(a_12_), .CI(n15), .CO(n14), .S(product_19_) );
  ADDFXL U20 ( .A(n158), .B(a_11_), .CI(n16), .CO(n15), .S(product_18_) );
  ADDFXL U21 ( .A(n32), .B(n163), .CI(n17), .CO(n16), .S(product_17_) );
  ADDFXL U22 ( .A(n34), .B(n33), .CI(n18), .CO(n17), .S(product_16_) );
  ADDFXL U23 ( .A(n35), .B(n36), .CI(n19), .CO(n18), .S(product_15_) );
  ADDFXL U24 ( .A(n37), .B(n38), .CI(n20), .CO(n19), .S(product_14_) );
  ADDFXL U25 ( .A(n39), .B(n40), .CI(n21), .CO(n20), .S(product_13_) );
  ADDFXL U26 ( .A(n41), .B(n42), .CI(n22), .CO(n21), .S(product_12_) );
  ADDFXL U27 ( .A(n43), .B(n44), .CI(n23), .CO(n22), .S(product_11_) );
  ADDFXL U28 ( .A(n45), .B(n46), .CI(n24), .CO(n23), .S(product_10_) );
  ADDFXL U29 ( .A(n47), .B(n48), .CI(n25), .CO(n24), .S(product_9_) );
  ADDFXL U30 ( .A(n49), .B(n50), .CI(n26), .CO(n25), .S(product_8_) );
  ADDFXL U31 ( .A(n51), .B(a_5_), .CI(n27), .CO(n26), .S(product_7_) );
  ADDFXL U32 ( .A(a_5_), .B(a_4_), .CI(n28), .CO(n27), .S(product_6_) );
  ADDFXL U33 ( .A(a_4_), .B(a_3_), .CI(n29), .CO(n28), .S(product_5_) );
  ADDFXL U34 ( .A(a_3_), .B(a_2_), .CI(n30), .CO(n29), .S(product_4_) );
  ADDFXL U35 ( .A(a_2_), .B(a_1_), .CI(n31), .CO(n30), .S(product_3_) );
  ADDHXL U36 ( .A(a_0_), .B(a_1_), .CO(n31), .S(product_2_) );
  ADDFXL U37 ( .A(n164), .B(a_15_), .CI(a_14_), .CO(n32), .S(n33) );
  ADDFXL U38 ( .A(a_13_), .B(n165), .CI(a_14_), .CO(n34), .S(n35) );
  ADDFXL U39 ( .A(a_12_), .B(n166), .CI(a_13_), .CO(n36), .S(n37) );
  ADDFXL U40 ( .A(a_11_), .B(n167), .CI(a_12_), .CO(n38), .S(n39) );
  ADDFXL U41 ( .A(a_10_), .B(n168), .CI(a_11_), .CO(n40), .S(n41) );
  ADDFXL U42 ( .A(a_9_), .B(n169), .CI(a_10_), .CO(n42), .S(n43) );
  ADDFXL U43 ( .A(a_8_), .B(n170), .CI(a_9_), .CO(n44), .S(n45) );
  ADDFXL U44 ( .A(a_7_), .B(n171), .CI(a_8_), .CO(n46), .S(n47) );
  ADDFXL U45 ( .A(a_6_), .B(n172), .CI(a_7_), .CO(n48), .S(n49) );
  INVX3 U68 ( .A(product_28_), .Y(n148) );
  CLKINVX1 U69 ( .A(n11), .Y(product_28_) );
  CLKINVX1 U70 ( .A(n148), .Y(product_23_) );
  CLKINVX1 U71 ( .A(n148), .Y(product_24_) );
  CLKINVX1 U72 ( .A(n148), .Y(product_25_) );
  CLKINVX1 U73 ( .A(n148), .Y(product_26_) );
  CLKINVX1 U74 ( .A(n148), .Y(product_27_) );
  CLKINVX1 U75 ( .A(n148), .Y(product_29_) );
  CLKINVX1 U76 ( .A(n148), .Y(product_30_) );
  CLKINVX1 U77 ( .A(n148), .Y(product_31_) );
  CLKINVX1 U78 ( .A(a_14_), .Y(n159) );
  CLKINVX1 U79 ( .A(a_13_), .Y(n160) );
  CLKINVX1 U80 ( .A(a_15_), .Y(n158) );
  CLKINVX1 U81 ( .A(a_11_), .Y(n162) );
  CLKINVX1 U82 ( .A(a_12_), .Y(n161) );
  CLKINVX1 U83 ( .A(a_10_), .Y(n163) );
  CLKINVX1 U84 ( .A(a_1_), .Y(n172) );
  CLKINVX1 U85 ( .A(a_2_), .Y(n171) );
  CLKINVX1 U86 ( .A(a_3_), .Y(n170) );
  CLKINVX1 U87 ( .A(a_4_), .Y(n169) );
  CLKINVX1 U88 ( .A(a_6_), .Y(n167) );
  CLKINVX1 U89 ( .A(a_5_), .Y(n168) );
  CLKINVX1 U90 ( .A(a_7_), .Y(n166) );
  CLKINVX1 U91 ( .A(a_9_), .Y(n164) );
  CLKINVX1 U92 ( .A(a_8_), .Y(n165) );
  CLKBUFX3 U93 ( .A(a_0_), .Y(product_1_) );
  XOR2X1 U94 ( .A(a_6_), .B(a_0_), .Y(n51) );
  NAND2X1 U95 ( .A(a_0_), .B(n167), .Y(n50) );
endmodule


module FIR_FILTER2_DW_mult_uns_13 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n176, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201;

  ADDFXL U16 ( .A(a_15_), .B(n187), .CI(n12), .CO(n11), .S(product_22_) );
  ADDFXL U17 ( .A(n34), .B(a_14_), .CI(n13), .CO(n12), .S(product_21_) );
  ADDFXL U18 ( .A(n35), .B(n36), .CI(n14), .CO(n13), .S(product_20_) );
  ADDFXL U19 ( .A(n37), .B(n39), .CI(n15), .CO(n14), .S(product_19_) );
  ADDFXL U20 ( .A(n40), .B(n42), .CI(n16), .CO(n15), .S(product_18_) );
  ADDFXL U21 ( .A(n43), .B(n45), .CI(n17), .CO(n16), .S(product_17_) );
  ADDFXL U22 ( .A(n46), .B(n48), .CI(n18), .CO(n17), .S(product_16_) );
  ADDFXL U23 ( .A(n49), .B(n51), .CI(n19), .CO(n18), .S(product_15_) );
  ADDFXL U24 ( .A(n52), .B(n54), .CI(n20), .CO(n19), .S(product_14_) );
  ADDFXL U25 ( .A(n55), .B(n57), .CI(n21), .CO(n20), .S(product_13_) );
  ADDFXL U26 ( .A(n58), .B(n60), .CI(n22), .CO(n21), .S(product_12_) );
  ADDFXL U27 ( .A(n61), .B(n63), .CI(n23), .CO(n22), .S(product_11_) );
  ADDFXL U28 ( .A(n64), .B(n66), .CI(n24), .CO(n23), .S(product_10_) );
  ADDFXL U29 ( .A(n67), .B(n69), .CI(n25), .CO(n24), .S(product_9_) );
  ADDFXL U30 ( .A(n71), .B(n70), .CI(n26), .CO(n25), .S(product_8_) );
  ADDFXL U31 ( .A(n72), .B(n75), .CI(n27), .CO(n26), .S(product_7_) );
  ADDFXL U32 ( .A(n76), .B(n77), .CI(n28), .CO(n27), .S(product_6_) );
  ADDFXL U33 ( .A(n78), .B(a_0_), .CI(n29), .CO(n28), .S(product_5_) );
  ADDFXL U34 ( .A(a_1_), .B(n197), .CI(n30), .CO(n29), .S(product_4_) );
  ADDFXL U35 ( .A(a_0_), .B(n198), .CI(n31), .CO(n30), .S(product_3_) );
  ADDHXL U36 ( .A(n199), .B(n32), .CO(n31), .S(product_2_) );
  ADDHXL U37 ( .A(n200), .B(n201), .CO(n32), .S(product_1_) );
  ADDFXL U39 ( .A(n189), .B(n186), .CI(n188), .CO(n34), .S(n35) );
  ADDFXL U40 ( .A(a_14_), .B(a_12_), .CI(n38), .CO(n36), .S(n37) );
  CMPR42X1 U41 ( .A(n190), .B(n191), .C(n186), .D(a_13_), .ICI(n41), .S(n40), 
        .ICO(n38), .CO(n39) );
  CMPR42X1 U42 ( .A(a_10_), .B(n192), .C(a_14_), .D(a_12_), .ICI(n44), .S(n43), 
        .ICO(n41), .CO(n42) );
  CMPR42X1 U43 ( .A(a_9_), .B(n193), .C(a_13_), .D(a_11_), .ICI(n47), .S(n46), 
        .ICO(n44), .CO(n45) );
  CMPR42X1 U44 ( .A(a_8_), .B(a_15_), .C(a_12_), .D(a_10_), .ICI(n50), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U45 ( .A(n187), .B(n194), .C(a_9_), .D(a_11_), .ICI(n53), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U46 ( .A(n188), .B(n195), .C(a_8_), .D(a_10_), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U47 ( .A(n189), .B(n196), .C(a_7_), .D(a_9_), .ICI(n59), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U48 ( .A(n190), .B(n197), .C(a_6_), .D(a_8_), .ICI(n62), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U49 ( .A(n191), .B(n198), .C(a_5_), .D(a_7_), .ICI(n65), .S(n64), 
        .ICO(n62), .CO(n63) );
  CMPR42X1 U50 ( .A(n192), .B(n199), .C(a_4_), .D(a_6_), .ICI(n68), .S(n67), 
        .ICO(n65), .CO(n66) );
  CMPR42X1 U51 ( .A(n193), .B(n200), .C(a_3_), .D(a_5_), .ICI(n73), .S(n70), 
        .ICO(n68), .CO(n69) );
  ADDFXL U52 ( .A(a_2_), .B(a_4_), .CI(n74), .CO(n71), .S(n72) );
  ADDFXL U55 ( .A(a_1_), .B(n195), .CI(a_3_), .CO(n75), .S(n76) );
  ADDHXL U56 ( .A(n196), .B(a_2_), .CO(n77), .S(n78) );
  INVX3 U77 ( .A(product_28_), .Y(n176) );
  CLKINVX1 U78 ( .A(n11), .Y(product_28_) );
  CLKINVX1 U79 ( .A(n176), .Y(product_23_) );
  CLKINVX1 U80 ( .A(n176), .Y(product_24_) );
  CLKINVX1 U81 ( .A(n176), .Y(product_25_) );
  CLKINVX1 U82 ( .A(n176), .Y(product_26_) );
  CLKINVX1 U83 ( .A(n176), .Y(product_27_) );
  CLKINVX1 U84 ( .A(n176), .Y(product_29_) );
  CLKINVX1 U85 ( .A(n176), .Y(product_30_) );
  CLKINVX1 U86 ( .A(n176), .Y(product_31_) );
  CLKINVX1 U87 ( .A(a_0_), .Y(n201) );
  CLKINVX1 U88 ( .A(a_3_), .Y(n198) );
  CLKINVX1 U89 ( .A(a_2_), .Y(n199) );
  CLKINVX1 U90 ( .A(a_1_), .Y(n200) );
  CLKINVX1 U91 ( .A(a_8_), .Y(n193) );
  CLKINVX1 U92 ( .A(a_7_), .Y(n194) );
  CLKINVX1 U93 ( .A(a_5_), .Y(n196) );
  CLKINVX1 U94 ( .A(a_6_), .Y(n195) );
  CLKINVX1 U95 ( .A(a_4_), .Y(n197) );
  CLKINVX1 U96 ( .A(a_9_), .Y(n192) );
  CLKINVX1 U97 ( .A(a_10_), .Y(n191) );
  CLKINVX1 U98 ( .A(a_11_), .Y(n190) );
  CLKINVX1 U99 ( .A(a_12_), .Y(n189) );
  CLKINVX1 U100 ( .A(a_14_), .Y(n187) );
  CLKINVX1 U101 ( .A(a_13_), .Y(n188) );
  CLKINVX1 U102 ( .A(a_15_), .Y(n186) );
  CLKBUFX3 U103 ( .A(a_0_), .Y(product_0_) );
  XOR2X1 U104 ( .A(n194), .B(a_0_), .Y(n74) );
  NAND2X1 U105 ( .A(a_0_), .B(a_7_), .Y(n73) );
endmodule


module FIR_FILTER2_DW_mult_uns_12 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n137, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  ADDFXL U17 ( .A(a_14_), .B(n148), .CI(n13), .CO(n12), .S(product_21_) );
  ADDFXL U18 ( .A(n149), .B(a_13_), .CI(n14), .CO(n13), .S(product_20_) );
  ADDFXL U19 ( .A(n150), .B(a_12_), .CI(n15), .CO(n14), .S(product_19_) );
  ADDFXL U20 ( .A(n40), .B(n151), .CI(n16), .CO(n15), .S(product_18_) );
  ADDFXL U21 ( .A(n41), .B(n42), .CI(n17), .CO(n16), .S(product_17_) );
  ADDFXL U22 ( .A(n44), .B(n43), .CI(n18), .CO(n17), .S(product_16_) );
  ADDFXL U23 ( .A(n46), .B(n45), .CI(n19), .CO(n18), .S(product_15_) );
  ADDFXL U24 ( .A(n47), .B(n48), .CI(n20), .CO(n19), .S(product_14_) );
  ADDFXL U25 ( .A(n49), .B(n50), .CI(n21), .CO(n20), .S(product_13_) );
  ADDFXL U26 ( .A(n51), .B(n52), .CI(n22), .CO(n21), .S(product_12_) );
  ADDFXL U27 ( .A(n53), .B(n54), .CI(n23), .CO(n22), .S(product_11_) );
  ADDFXL U28 ( .A(n55), .B(n56), .CI(n24), .CO(n23), .S(product_10_) );
  ADDFXL U29 ( .A(n57), .B(n58), .CI(n25), .CO(n24), .S(product_9_) );
  ADDFXL U30 ( .A(n59), .B(n60), .CI(n26), .CO(n25), .S(product_8_) );
  ADDFXL U31 ( .A(n61), .B(n62), .CI(n27), .CO(n26), .S(product_7_) );
  ADDFXL U32 ( .A(n63), .B(n64), .CI(n28), .CO(n27), .S(product_6_) );
  ADDFXL U33 ( .A(n65), .B(n66), .CI(n29), .CO(n28), .S(product_5_) );
  ADDFXL U34 ( .A(n67), .B(n68), .CI(n30), .CO(n29), .S(product_4_) );
  ADDFXL U35 ( .A(n69), .B(n161), .CI(n31), .CO(n30), .S(product_3_) );
  ADDFXL U36 ( .A(n163), .B(a_2_), .CI(n32), .CO(n31), .S(product_2_) );
  ADDHXL U37 ( .A(n162), .B(n163), .CO(n32), .S(product_1_) );
  ADDFXL U42 ( .A(a_11_), .B(n149), .CI(a_15_), .CO(n40), .S(n41) );
  ADDFXL U43 ( .A(n150), .B(a_14_), .CI(a_10_), .CO(n42), .S(n43) );
  ADDFXL U44 ( .A(a_9_), .B(a_13_), .CI(a_15_), .CO(n44), .S(n45) );
  ADDFXL U45 ( .A(n151), .B(n149), .CI(a_8_), .CO(n46), .S(n47) );
  ADDFXL U46 ( .A(n152), .B(n150), .CI(a_7_), .CO(n48), .S(n49) );
  ADDFXL U47 ( .A(n153), .B(n151), .CI(a_6_), .CO(n50), .S(n51) );
  ADDFXL U48 ( .A(n154), .B(n152), .CI(a_5_), .CO(n52), .S(n53) );
  ADDFXL U49 ( .A(n155), .B(n153), .CI(a_4_), .CO(n54), .S(n55) );
  ADDFXL U50 ( .A(n156), .B(n154), .CI(a_3_), .CO(n56), .S(n57) );
  ADDFXL U51 ( .A(n157), .B(n155), .CI(a_2_), .CO(n58), .S(n59) );
  ADDFXL U52 ( .A(n158), .B(n156), .CI(a_1_), .CO(n60), .S(n61) );
  ADDFXL U53 ( .A(n159), .B(n157), .CI(a_0_), .CO(n62), .S(n63) );
  ADDHXL U54 ( .A(n158), .B(n160), .CO(n64), .S(n65) );
  ADDHXL U55 ( .A(n159), .B(n161), .CO(n66), .S(n67) );
  ADDHXL U56 ( .A(n160), .B(n162), .CO(n68), .S(n69) );
  INVX3 U77 ( .A(product_29_), .Y(n137) );
  CLKINVX1 U78 ( .A(n137), .Y(product_22_) );
  CLKINVX1 U79 ( .A(n137), .Y(product_23_) );
  CLKINVX1 U80 ( .A(n137), .Y(product_24_) );
  CLKINVX1 U81 ( .A(n137), .Y(product_25_) );
  CLKINVX1 U82 ( .A(n137), .Y(product_26_) );
  CLKINVX1 U83 ( .A(n137), .Y(product_27_) );
  CLKINVX1 U84 ( .A(n137), .Y(product_28_) );
  CLKINVX1 U85 ( .A(n137), .Y(product_30_) );
  CLKINVX1 U86 ( .A(n137), .Y(product_31_) );
  CLKINVX1 U87 ( .A(n12), .Y(product_29_) );
  CLKINVX1 U88 ( .A(a_15_), .Y(n148) );
  CLKINVX1 U89 ( .A(a_0_), .Y(n163) );
  CLKINVX1 U90 ( .A(a_1_), .Y(n162) );
  CLKINVX1 U91 ( .A(a_2_), .Y(n161) );
  CLKINVX1 U92 ( .A(a_3_), .Y(n160) );
  CLKINVX1 U93 ( .A(a_4_), .Y(n159) );
  CLKINVX1 U94 ( .A(a_5_), .Y(n158) );
  CLKINVX1 U95 ( .A(a_6_), .Y(n157) );
  CLKINVX1 U96 ( .A(a_7_), .Y(n156) );
  CLKINVX1 U97 ( .A(a_8_), .Y(n155) );
  CLKINVX1 U98 ( .A(a_10_), .Y(n153) );
  CLKINVX1 U99 ( .A(a_9_), .Y(n154) );
  CLKINVX1 U100 ( .A(a_13_), .Y(n150) );
  CLKINVX1 U101 ( .A(a_12_), .Y(n151) );
  CLKINVX1 U102 ( .A(a_11_), .Y(n152) );
  CLKINVX1 U103 ( .A(a_14_), .Y(n149) );
  CLKBUFX3 U104 ( .A(a_0_), .Y(product_0_) );
endmodule


module FIR_FILTER2_DW_mult_uns_11 ( a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_,
         a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n172;

  ADDFXL U16 ( .A(a_14_), .B(a_15_), .CI(n12), .CO(product_23_), .S(
        product_22_) );
  ADDFXL U17 ( .A(n33), .B(a_13_), .CI(n13), .CO(n12), .S(product_21_) );
  ADDFXL U18 ( .A(n35), .B(n34), .CI(n14), .CO(n13), .S(product_20_) );
  ADDFXL U19 ( .A(n37), .B(n36), .CI(n15), .CO(n14), .S(product_19_) );
  ADDFXL U20 ( .A(n38), .B(n40), .CI(n16), .CO(n15), .S(product_18_) );
  ADDFXL U21 ( .A(n43), .B(n41), .CI(n17), .CO(n16), .S(product_17_) );
  ADDFXL U22 ( .A(n44), .B(n46), .CI(n18), .CO(n17), .S(product_16_) );
  ADDFXL U23 ( .A(n47), .B(n51), .CI(n19), .CO(n18), .S(product_15_) );
  ADDFXL U24 ( .A(n52), .B(n56), .CI(n20), .CO(n19), .S(product_14_) );
  ADDFXL U25 ( .A(n57), .B(n61), .CI(n21), .CO(n20), .S(product_13_) );
  ADDFXL U26 ( .A(n62), .B(n66), .CI(n22), .CO(n21), .S(product_12_) );
  ADDFXL U27 ( .A(n67), .B(n71), .CI(n23), .CO(n22), .S(product_11_) );
  ADDFXL U28 ( .A(n72), .B(n76), .CI(n24), .CO(n23), .S(product_10_) );
  ADDFXL U29 ( .A(n77), .B(n81), .CI(n25), .CO(n24), .S(product_9_) );
  ADDFXL U30 ( .A(n82), .B(n86), .CI(n26), .CO(n25), .S(product_8_) );
  ADDFXL U31 ( .A(n88), .B(n87), .CI(n27), .CO(n26), .S(product_7_) );
  ADDFXL U32 ( .A(n89), .B(n92), .CI(n28), .CO(n27), .S(product_6_) );
  ADDFXL U33 ( .A(n93), .B(n94), .CI(n29), .CO(n28), .S(product_5_) );
  ADDFXL U34 ( .A(n95), .B(n96), .CI(n30), .CO(n29), .S(product_4_) );
  ADDFXL U35 ( .A(n97), .B(a_0_), .CI(n31), .CO(n30), .S(product_3_) );
  ADDFXL U36 ( .A(a_2_), .B(a_1_), .CI(n32), .CO(n31), .S(product_2_) );
  ADDHXL U37 ( .A(a_0_), .B(a_1_), .CO(n32), .S(product_1_) );
  ADDFXL U38 ( .A(a_14_), .B(a_15_), .CI(a_12_), .CO(n33), .S(n34) );
  ADDFXL U39 ( .A(a_13_), .B(a_15_), .CI(a_11_), .CO(n35), .S(n36) );
  ADDFXL U40 ( .A(a_10_), .B(a_12_), .CI(n39), .CO(n37), .S(n38) );
  CMPR42X1 U41 ( .A(a_15_), .B(a_14_), .C(a_9_), .D(a_11_), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U42 ( .A(a_13_), .B(a_8_), .C(a_10_), .D(n48), .ICI(n45), .S(n44), 
        .ICO(n42), .CO(n43) );
  CMPR42X1 U43 ( .A(a_14_), .B(a_12_), .C(n49), .D(n53), .ICI(n50), .S(n47), 
        .ICO(n45), .CO(n46) );
  ADDFXL U44 ( .A(a_9_), .B(a_15_), .CI(a_7_), .CO(n48), .S(n49) );
  CMPR42X1 U45 ( .A(a_14_), .B(a_13_), .C(n58), .D(n54), .ICI(n55), .S(n52), 
        .ICO(n50), .CO(n51) );
  ADDFXL U46 ( .A(a_6_), .B(a_8_), .CI(a_11_), .CO(n53), .S(n54) );
  CMPR42X1 U47 ( .A(a_13_), .B(a_12_), .C(n63), .D(n59), .ICI(n60), .S(n57), 
        .ICO(n55), .CO(n56) );
  ADDFXL U48 ( .A(a_5_), .B(a_7_), .CI(a_10_), .CO(n58), .S(n59) );
  CMPR42X1 U49 ( .A(a_12_), .B(a_11_), .C(n68), .D(n64), .ICI(n65), .S(n62), 
        .ICO(n60), .CO(n61) );
  ADDFXL U50 ( .A(a_4_), .B(a_6_), .CI(a_9_), .CO(n63), .S(n64) );
  CMPR42X1 U51 ( .A(a_11_), .B(a_10_), .C(n73), .D(n69), .ICI(n70), .S(n67), 
        .ICO(n65), .CO(n66) );
  ADDFXL U52 ( .A(a_3_), .B(a_5_), .CI(a_8_), .CO(n68), .S(n69) );
  CMPR42X1 U53 ( .A(a_10_), .B(a_9_), .C(n75), .D(n78), .ICI(n74), .S(n72), 
        .ICO(n70), .CO(n71) );
  ADDFXL U54 ( .A(a_2_), .B(a_4_), .CI(a_7_), .CO(n73), .S(n74) );
  CMPR42X1 U55 ( .A(a_9_), .B(a_8_), .C(n83), .D(n80), .ICI(n79), .S(n77), 
        .ICO(n75), .CO(n76) );
  ADDFXL U56 ( .A(a_1_), .B(a_3_), .CI(a_6_), .CO(n78), .S(n79) );
  CMPR42X1 U57 ( .A(a_8_), .B(a_5_), .C(a_7_), .D(n85), .ICI(n84), .S(n82), 
        .ICO(n80), .CO(n81) );
  ADDHXL U58 ( .A(a_2_), .B(a_0_), .CO(n83), .S(n84) );
  CMPR42X1 U59 ( .A(a_4_), .B(a_1_), .C(a_6_), .D(a_7_), .ICI(n90), .S(n87), 
        .ICO(n85), .CO(n86) );
  ADDFXL U60 ( .A(a_5_), .B(a_6_), .CI(n91), .CO(n88), .S(n89) );
  ADDHXL U61 ( .A(a_3_), .B(a_0_), .CO(n90), .S(n91) );
  ADDFXL U62 ( .A(a_2_), .B(a_5_), .CI(a_4_), .CO(n92), .S(n93) );
  ADDFXL U63 ( .A(a_1_), .B(a_4_), .CI(a_3_), .CO(n94), .S(n95) );
  ADDHXL U64 ( .A(a_3_), .B(a_2_), .CO(n96), .S(n97) );
  INVX3 U85 ( .A(a_16_), .Y(n172) );
  CLKINVX1 U86 ( .A(n172), .Y(product_24_) );
  CLKINVX1 U87 ( .A(n172), .Y(product_25_) );
  CLKINVX1 U88 ( .A(n172), .Y(product_26_) );
  CLKINVX1 U89 ( .A(n172), .Y(product_27_) );
  CLKINVX1 U90 ( .A(n172), .Y(product_28_) );
  CLKINVX1 U91 ( .A(n172), .Y(product_29_) );
  CLKINVX1 U92 ( .A(n172), .Y(product_30_) );
  CLKINVX1 U93 ( .A(n172), .Y(product_31_) );
  CLKBUFX3 U94 ( .A(a_0_), .Y(product_0_) );
endmodule


module FIR_FILTER2_DW_mult_uns_10 ( a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_,
         a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n126;

  ADDFXL U11 ( .A(a_14_), .B(a_15_), .CI(n9), .CO(product_24_), .S(product_23_) );
  ADDFXL U12 ( .A(a_13_), .B(a_15_), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U13 ( .A(n29), .B(a_12_), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U14 ( .A(n31), .B(n30), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U15 ( .A(n33), .B(n32), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U16 ( .A(n34), .B(n36), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U17 ( .A(n37), .B(n39), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U18 ( .A(n42), .B(n40), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U19 ( .A(n43), .B(n45), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U20 ( .A(n46), .B(n48), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U21 ( .A(n49), .B(n51), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U22 ( .A(n52), .B(n54), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U23 ( .A(n55), .B(n57), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U24 ( .A(n59), .B(n58), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U25 ( .A(n60), .B(n63), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U26 ( .A(n64), .B(n65), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U27 ( .A(n66), .B(n67), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U28 ( .A(n68), .B(a_0_), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFXL U29 ( .A(a_4_), .B(a_2_), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFXL U30 ( .A(a_3_), .B(a_1_), .CI(n28), .CO(n27), .S(product_4_) );
  ADDHXL U31 ( .A(a_0_), .B(a_2_), .CO(n28), .S(product_3_) );
  ADDFXL U32 ( .A(a_14_), .B(a_15_), .CI(a_11_), .CO(n29), .S(n30) );
  ADDFXL U33 ( .A(a_13_), .B(a_15_), .CI(a_10_), .CO(n31), .S(n32) );
  ADDFXL U34 ( .A(a_9_), .B(a_12_), .CI(n35), .CO(n33), .S(n34) );
  CMPR42X1 U35 ( .A(a_15_), .B(a_14_), .C(a_8_), .D(a_11_), .ICI(n38), .S(n37), 
        .ICO(n35), .CO(n36) );
  CMPR42X1 U36 ( .A(a_15_), .B(a_13_), .C(a_7_), .D(a_10_), .ICI(n41), .S(n40), 
        .ICO(n38), .CO(n39) );
  CMPR42X1 U37 ( .A(a_9_), .B(a_6_), .C(a_12_), .D(a_14_), .ICI(n44), .S(n43), 
        .ICO(n41), .CO(n42) );
  CMPR42X1 U38 ( .A(a_8_), .B(a_5_), .C(a_11_), .D(a_13_), .ICI(n47), .S(n46), 
        .ICO(n44), .CO(n45) );
  CMPR42X1 U39 ( .A(a_7_), .B(a_4_), .C(a_10_), .D(a_12_), .ICI(n50), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U40 ( .A(a_6_), .B(a_3_), .C(a_9_), .D(a_11_), .ICI(n53), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U41 ( .A(a_5_), .B(a_2_), .C(a_8_), .D(a_10_), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U42 ( .A(a_4_), .B(a_1_), .C(a_7_), .D(a_9_), .ICI(n61), .S(n58), 
        .ICO(n56), .CO(n57) );
  ADDFXL U43 ( .A(a_6_), .B(a_8_), .CI(n62), .CO(n59), .S(n60) );
  ADDHXL U44 ( .A(a_3_), .B(a_0_), .CO(n61), .S(n62) );
  ADDFXL U45 ( .A(a_2_), .B(a_7_), .CI(a_5_), .CO(n63), .S(n64) );
  ADDFXL U46 ( .A(a_1_), .B(a_6_), .CI(a_4_), .CO(n65), .S(n66) );
  ADDHXL U47 ( .A(a_5_), .B(a_3_), .CO(n67), .S(n68) );
  INVX3 U53 ( .A(a_16_), .Y(n126) );
  CLKINVX1 U54 ( .A(n126), .Y(product_25_) );
  CLKINVX1 U55 ( .A(n126), .Y(product_26_) );
  CLKINVX1 U56 ( .A(n126), .Y(product_27_) );
  CLKINVX1 U57 ( .A(n126), .Y(product_28_) );
  CLKINVX1 U58 ( .A(n126), .Y(product_29_) );
  CLKINVX1 U59 ( .A(n126), .Y(product_30_) );
  CLKINVX1 U60 ( .A(n126), .Y(product_31_) );
  CLKBUFX3 U61 ( .A(a_1_), .Y(product_2_) );
  CLKBUFX3 U62 ( .A(a_0_), .Y(product_1_) );
endmodule


module FIR_FILTER2_DW_mult_uns_9 ( a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_,
         a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n104;

  ADDFXL U11 ( .A(a_14_), .B(a_15_), .CI(n9), .CO(product_24_), .S(product_23_) );
  ADDFXL U12 ( .A(a_13_), .B(a_15_), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U13 ( .A(a_12_), .B(a_15_), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U14 ( .A(n27), .B(a_11_), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U15 ( .A(n29), .B(n28), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U16 ( .A(n31), .B(n30), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U17 ( .A(n33), .B(n32), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U18 ( .A(n35), .B(n34), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U19 ( .A(n36), .B(n37), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U20 ( .A(n38), .B(n39), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U21 ( .A(n40), .B(n41), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U22 ( .A(n42), .B(n43), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U23 ( .A(n44), .B(n45), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U24 ( .A(n46), .B(n47), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U25 ( .A(n48), .B(a_0_), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U26 ( .A(a_7_), .B(a_3_), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U27 ( .A(a_6_), .B(a_2_), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U28 ( .A(a_5_), .B(a_1_), .CI(n26), .CO(n25), .S(product_6_) );
  ADDHXL U29 ( .A(a_0_), .B(a_4_), .CO(n26), .S(product_5_) );
  ADDFXL U30 ( .A(a_14_), .B(a_15_), .CI(a_10_), .CO(n27), .S(n28) );
  ADDFXL U31 ( .A(a_13_), .B(a_15_), .CI(a_9_), .CO(n29), .S(n30) );
  ADDFXL U32 ( .A(a_12_), .B(a_15_), .CI(a_8_), .CO(n31), .S(n32) );
  ADDFXL U33 ( .A(a_11_), .B(a_15_), .CI(a_7_), .CO(n33), .S(n34) );
  ADDFXL U34 ( .A(a_6_), .B(a_14_), .CI(a_10_), .CO(n35), .S(n36) );
  ADDFXL U35 ( .A(a_5_), .B(a_13_), .CI(a_9_), .CO(n37), .S(n38) );
  ADDFXL U36 ( .A(a_4_), .B(a_12_), .CI(a_8_), .CO(n39), .S(n40) );
  ADDFXL U37 ( .A(a_3_), .B(a_11_), .CI(a_7_), .CO(n41), .S(n42) );
  ADDFXL U38 ( .A(a_2_), .B(a_10_), .CI(a_6_), .CO(n43), .S(n44) );
  ADDFXL U39 ( .A(a_1_), .B(a_9_), .CI(a_5_), .CO(n45), .S(n46) );
  ADDHXL U40 ( .A(a_8_), .B(a_4_), .CO(n47), .S(n48) );
  INVX3 U46 ( .A(a_16_), .Y(n104) );
  CLKINVX1 U47 ( .A(n104), .Y(product_25_) );
  CLKINVX1 U48 ( .A(n104), .Y(product_26_) );
  CLKINVX1 U49 ( .A(n104), .Y(product_27_) );
  CLKINVX1 U50 ( .A(n104), .Y(product_28_) );
  CLKINVX1 U51 ( .A(n104), .Y(product_29_) );
  CLKINVX1 U52 ( .A(n104), .Y(product_30_) );
  CLKINVX1 U53 ( .A(n104), .Y(product_31_) );
  CLKBUFX3 U54 ( .A(a_3_), .Y(product_4_) );
  CLKBUFX3 U55 ( .A(a_2_), .Y(product_3_) );
  CLKBUFX3 U56 ( .A(a_1_), .Y(product_2_) );
  CLKBUFX3 U57 ( .A(a_0_), .Y(product_1_) );
endmodule


module FIR_FILTER2_DW_mult_uns_7 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n173, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195;

  ADDFXL U11 ( .A(a_15_), .B(n182), .CI(n8), .CO(n7), .S(product_25_) );
  ADDFXL U12 ( .A(n183), .B(a_14_), .CI(n9), .CO(n8), .S(product_24_) );
  ADDFXL U13 ( .A(n184), .B(a_13_), .CI(n10), .CO(n9), .S(product_23_) );
  ADDFXL U14 ( .A(n31), .B(a_12_), .CI(n11), .CO(n10), .S(product_22_) );
  ADDFXL U15 ( .A(n32), .B(n33), .CI(n12), .CO(n11), .S(product_21_) );
  ADDFXL U16 ( .A(n35), .B(n34), .CI(n13), .CO(n12), .S(product_20_) );
  ADDFXL U17 ( .A(n37), .B(n36), .CI(n14), .CO(n13), .S(product_19_) );
  ADDFXL U18 ( .A(n38), .B(n40), .CI(n15), .CO(n14), .S(product_18_) );
  ADDFXL U19 ( .A(n41), .B(n43), .CI(n16), .CO(n15), .S(product_17_) );
  ADDFXL U20 ( .A(n44), .B(n46), .CI(n17), .CO(n16), .S(product_16_) );
  ADDFXL U21 ( .A(n49), .B(n47), .CI(n18), .CO(n17), .S(product_15_) );
  ADDFXL U22 ( .A(n50), .B(n52), .CI(n19), .CO(n18), .S(product_14_) );
  ADDFXL U23 ( .A(n53), .B(n55), .CI(n20), .CO(n19), .S(product_13_) );
  ADDFXL U24 ( .A(n56), .B(n58), .CI(n21), .CO(n20), .S(product_12_) );
  ADDFXL U25 ( .A(n60), .B(n59), .CI(n22), .CO(n21), .S(product_11_) );
  ADDFXL U26 ( .A(n61), .B(n64), .CI(n23), .CO(n22), .S(product_10_) );
  ADDFXL U27 ( .A(n65), .B(n66), .CI(n24), .CO(n23), .S(product_9_) );
  ADDFXL U28 ( .A(n67), .B(n68), .CI(n25), .CO(n24), .S(product_8_) );
  ADDFXL U29 ( .A(n69), .B(n70), .CI(n26), .CO(n25), .S(product_7_) );
  ADDFXL U30 ( .A(n71), .B(a_4_), .CI(n27), .CO(n26), .S(product_6_) );
  ADDFXL U31 ( .A(a_5_), .B(a_3_), .CI(n28), .CO(n27), .S(product_5_) );
  ADDFXL U32 ( .A(a_4_), .B(a_2_), .CI(n29), .CO(n28), .S(product_4_) );
  ADDFXL U33 ( .A(a_3_), .B(a_1_), .CI(n30), .CO(n29), .S(product_3_) );
  ADDHXL U34 ( .A(a_0_), .B(a_2_), .CO(n30), .S(product_2_) );
  ADDFXL U35 ( .A(n185), .B(n182), .CI(a_15_), .CO(n31), .S(n32) );
  ADDFXL U36 ( .A(n186), .B(a_14_), .CI(n183), .CO(n33), .S(n34) );
  ADDFXL U37 ( .A(n187), .B(a_13_), .CI(n184), .CO(n35), .S(n36) );
  ADDFXL U38 ( .A(n188), .B(a_12_), .CI(n39), .CO(n37), .S(n38) );
  CMPR42X1 U39 ( .A(n189), .B(n186), .C(n185), .D(n181), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U40 ( .A(a_10_), .B(n181), .C(n190), .D(a_14_), .ICI(n45), .S(n44), 
        .ICO(n42), .CO(n43) );
  CMPR42X1 U41 ( .A(a_15_), .B(n191), .C(n187), .D(a_13_), .ICI(n48), .S(n47), 
        .ICO(n45), .CO(n46) );
  CMPR42X1 U42 ( .A(n192), .B(n188), .C(a_12_), .D(a_14_), .ICI(n51), .S(n50), 
        .ICO(n48), .CO(n49) );
  CMPR42X1 U43 ( .A(n193), .B(n189), .C(a_11_), .D(a_13_), .ICI(n54), .S(n53), 
        .ICO(n51), .CO(n52) );
  CMPR42X1 U44 ( .A(n194), .B(n190), .C(a_10_), .D(a_12_), .ICI(n57), .S(n56), 
        .ICO(n54), .CO(n55) );
  CMPR42X1 U45 ( .A(n195), .B(n191), .C(a_9_), .D(a_11_), .ICI(n62), .S(n59), 
        .ICO(n57), .CO(n58) );
  ADDFXL U46 ( .A(a_8_), .B(a_10_), .CI(n63), .CO(n60), .S(n61) );
  ADDFXL U49 ( .A(a_7_), .B(n193), .CI(a_9_), .CO(n64), .S(n65) );
  ADDFXL U50 ( .A(a_6_), .B(n194), .CI(a_8_), .CO(n66), .S(n67) );
  ADDFXL U51 ( .A(a_5_), .B(n195), .CI(a_7_), .CO(n68), .S(n69) );
  CLKINVX1 U77 ( .A(product_28_), .Y(n173) );
  CLKINVX1 U78 ( .A(n173), .Y(product_26_) );
  CLKINVX1 U79 ( .A(n173), .Y(product_27_) );
  CLKINVX1 U80 ( .A(n173), .Y(product_29_) );
  CLKINVX1 U81 ( .A(n173), .Y(product_30_) );
  CLKINVX1 U82 ( .A(n173), .Y(product_31_) );
  CLKINVX1 U83 ( .A(a_6_), .Y(n190) );
  CLKINVX1 U84 ( .A(a_2_), .Y(n194) );
  CLKINVX1 U85 ( .A(a_1_), .Y(n195) );
  CLKINVX1 U86 ( .A(a_5_), .Y(n191) );
  CLKINVX1 U87 ( .A(a_4_), .Y(n192) );
  CLKINVX1 U88 ( .A(a_3_), .Y(n193) );
  CLKINVX1 U89 ( .A(a_7_), .Y(n189) );
  CLKINVX1 U90 ( .A(a_8_), .Y(n188) );
  CLKINVX1 U91 ( .A(a_15_), .Y(n181) );
  CLKINVX1 U92 ( .A(a_10_), .Y(n186) );
  CLKINVX1 U93 ( .A(a_11_), .Y(n185) );
  CLKINVX1 U94 ( .A(a_9_), .Y(n187) );
  CLKINVX1 U95 ( .A(a_12_), .Y(n184) );
  CLKINVX1 U96 ( .A(a_13_), .Y(n183) );
  CLKINVX1 U97 ( .A(a_14_), .Y(n182) );
  CLKBUFX3 U98 ( .A(a_1_), .Y(product_1_) );
  CLKBUFX3 U99 ( .A(a_0_), .Y(product_0_) );
  CLKINVX1 U100 ( .A(n7), .Y(product_28_) );
  XOR2X1 U101 ( .A(a_6_), .B(a_0_), .Y(n71) );
  NAND2X1 U102 ( .A(a_0_), .B(n190), .Y(n70) );
  XOR2X1 U103 ( .A(n192), .B(a_0_), .Y(n63) );
  NAND2X1 U104 ( .A(a_0_), .B(a_4_), .Y(n62) );
endmodule


module FIR_FILTER2_DW_mult_uns_6 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n171, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192;

  ADDFXL U9 ( .A(a_15_), .B(n179), .CI(n7), .CO(n6), .S(product_26_) );
  ADDFXL U10 ( .A(n180), .B(a_14_), .CI(n8), .CO(n7), .S(product_25_) );
  ADDFXL U11 ( .A(n181), .B(a_13_), .CI(n9), .CO(n8), .S(product_24_) );
  ADDFXL U12 ( .A(n182), .B(a_12_), .CI(n10), .CO(n9), .S(product_23_) );
  ADDFXL U13 ( .A(n30), .B(a_11_), .CI(n11), .CO(n10), .S(product_22_) );
  ADDFXL U14 ( .A(n31), .B(n32), .CI(n12), .CO(n11), .S(product_21_) );
  ADDFXL U15 ( .A(n34), .B(n33), .CI(n13), .CO(n12), .S(product_20_) );
  ADDFXL U16 ( .A(n35), .B(n37), .CI(n14), .CO(n13), .S(product_19_) );
  ADDFXL U17 ( .A(n38), .B(n40), .CI(n15), .CO(n14), .S(product_18_) );
  ADDFXL U18 ( .A(n41), .B(n43), .CI(n16), .CO(n15), .S(product_17_) );
  ADDFXL U19 ( .A(n46), .B(n44), .CI(n17), .CO(n16), .S(product_16_) );
  ADDFXL U20 ( .A(n47), .B(n49), .CI(n18), .CO(n17), .S(product_15_) );
  ADDFXL U21 ( .A(n50), .B(n52), .CI(n19), .CO(n18), .S(product_14_) );
  ADDFXL U22 ( .A(n53), .B(n55), .CI(n20), .CO(n19), .S(product_13_) );
  ADDFXL U23 ( .A(n57), .B(n56), .CI(n21), .CO(n20), .S(product_12_) );
  ADDFXL U24 ( .A(n58), .B(n61), .CI(n22), .CO(n21), .S(product_11_) );
  ADDFXL U25 ( .A(n62), .B(n63), .CI(n23), .CO(n22), .S(product_10_) );
  ADDFXL U26 ( .A(n64), .B(n65), .CI(n24), .CO(n23), .S(product_9_) );
  ADDFXL U27 ( .A(n66), .B(n67), .CI(n25), .CO(n24), .S(product_8_) );
  ADDFXL U28 ( .A(n68), .B(n69), .CI(n26), .CO(n25), .S(product_7_) );
  ADDFXL U29 ( .A(n70), .B(a_3_), .CI(n27), .CO(n26), .S(product_6_) );
  ADDFXL U30 ( .A(a_4_), .B(a_2_), .CI(n28), .CO(n27), .S(product_5_) );
  ADDFXL U31 ( .A(a_3_), .B(a_1_), .CI(n29), .CO(n28), .S(product_4_) );
  ADDHXL U32 ( .A(a_0_), .B(a_2_), .CO(n29), .S(product_3_) );
  ADDFXL U33 ( .A(n183), .B(n179), .CI(a_15_), .CO(n30), .S(n31) );
  ADDFXL U34 ( .A(n184), .B(a_14_), .CI(n180), .CO(n32), .S(n33) );
  ADDFXL U35 ( .A(n185), .B(a_13_), .CI(n36), .CO(n34), .S(n35) );
  CMPR42X1 U36 ( .A(n186), .B(n182), .C(n181), .D(n178), .ICI(n39), .S(n38), 
        .ICO(n36), .CO(n37) );
  CMPR42X1 U37 ( .A(a_11_), .B(n178), .C(n187), .D(a_14_), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U38 ( .A(a_15_), .B(n188), .C(n183), .D(a_13_), .ICI(n45), .S(n44), 
        .ICO(n42), .CO(n43) );
  CMPR42X1 U39 ( .A(n189), .B(n184), .C(a_12_), .D(a_14_), .ICI(n48), .S(n47), 
        .ICO(n45), .CO(n46) );
  CMPR42X1 U40 ( .A(n190), .B(n185), .C(a_11_), .D(a_13_), .ICI(n51), .S(n50), 
        .ICO(n48), .CO(n49) );
  CMPR42X1 U41 ( .A(n191), .B(n186), .C(a_10_), .D(a_12_), .ICI(n54), .S(n53), 
        .ICO(n51), .CO(n52) );
  CMPR42X1 U42 ( .A(n192), .B(n187), .C(a_9_), .D(a_11_), .ICI(n59), .S(n56), 
        .ICO(n54), .CO(n55) );
  ADDFXL U43 ( .A(a_8_), .B(a_10_), .CI(n60), .CO(n57), .S(n58) );
  ADDFXL U46 ( .A(a_7_), .B(n189), .CI(a_9_), .CO(n61), .S(n62) );
  ADDFXL U47 ( .A(a_6_), .B(n190), .CI(a_8_), .CO(n63), .S(n64) );
  ADDFXL U48 ( .A(a_5_), .B(n191), .CI(a_7_), .CO(n65), .S(n66) );
  ADDFXL U49 ( .A(a_4_), .B(n192), .CI(a_6_), .CO(n67), .S(n68) );
  CLKINVX1 U75 ( .A(product_28_), .Y(n171) );
  CLKINVX1 U76 ( .A(n171), .Y(product_27_) );
  CLKINVX1 U77 ( .A(n171), .Y(product_29_) );
  CLKINVX1 U78 ( .A(n171), .Y(product_30_) );
  CLKINVX1 U79 ( .A(n171), .Y(product_31_) );
  CLKINVX1 U80 ( .A(a_5_), .Y(n188) );
  CLKINVX1 U81 ( .A(a_2_), .Y(n191) );
  CLKINVX1 U82 ( .A(a_1_), .Y(n192) );
  CLKINVX1 U83 ( .A(a_3_), .Y(n190) );
  CLKINVX1 U84 ( .A(a_6_), .Y(n187) );
  CLKINVX1 U85 ( .A(a_4_), .Y(n189) );
  CLKINVX1 U86 ( .A(a_7_), .Y(n186) );
  CLKINVX1 U87 ( .A(a_9_), .Y(n184) );
  CLKINVX1 U88 ( .A(a_8_), .Y(n185) );
  CLKINVX1 U89 ( .A(a_11_), .Y(n182) );
  CLKINVX1 U90 ( .A(a_15_), .Y(n178) );
  CLKINVX1 U91 ( .A(a_12_), .Y(n181) );
  CLKINVX1 U92 ( .A(a_10_), .Y(n183) );
  CLKINVX1 U93 ( .A(a_13_), .Y(n180) );
  CLKINVX1 U94 ( .A(a_14_), .Y(n179) );
  CLKBUFX3 U95 ( .A(a_1_), .Y(product_2_) );
  CLKBUFX3 U96 ( .A(a_0_), .Y(product_1_) );
  CLKINVX1 U97 ( .A(n6), .Y(product_28_) );
  XNOR2X1 U98 ( .A(n188), .B(a_0_), .Y(n70) );
  NAND2X1 U99 ( .A(a_0_), .B(n188), .Y(n69) );
  XNOR2X1 U100 ( .A(a_0_), .B(a_5_), .Y(n60) );
  NAND2X1 U101 ( .A(a_0_), .B(a_5_), .Y(n59) );
endmodule


module FIR_FILTER2_DW_mult_uns_5 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n201, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222;

  ADDFXL U9 ( .A(a_15_), .B(n208), .CI(n7), .CO(n6), .S(product_26_) );
  ADDFXL U10 ( .A(n209), .B(a_14_), .CI(n8), .CO(n7), .S(product_25_) );
  ADDFXL U11 ( .A(n32), .B(a_13_), .CI(n9), .CO(n8), .S(product_24_) );
  ADDFXL U12 ( .A(n33), .B(n34), .CI(n10), .CO(n9), .S(product_23_) );
  ADDFXL U13 ( .A(n35), .B(n37), .CI(n11), .CO(n10), .S(product_22_) );
  ADDFXL U14 ( .A(n40), .B(n38), .CI(n12), .CO(n11), .S(product_21_) );
  ADDFXL U15 ( .A(n41), .B(n43), .CI(n13), .CO(n12), .S(product_20_) );
  ADDFXL U16 ( .A(n44), .B(n48), .CI(n14), .CO(n13), .S(product_19_) );
  ADDFXL U17 ( .A(n49), .B(n53), .CI(n15), .CO(n14), .S(product_18_) );
  ADDFXL U18 ( .A(n54), .B(n58), .CI(n16), .CO(n15), .S(product_17_) );
  ADDFXL U19 ( .A(n59), .B(n63), .CI(n17), .CO(n16), .S(product_16_) );
  ADDFXL U20 ( .A(n64), .B(n68), .CI(n18), .CO(n17), .S(product_15_) );
  ADDFXL U21 ( .A(n69), .B(n73), .CI(n19), .CO(n18), .S(product_14_) );
  ADDFXL U22 ( .A(n74), .B(n78), .CI(n20), .CO(n19), .S(product_13_) );
  ADDFXL U23 ( .A(n79), .B(n83), .CI(n21), .CO(n20), .S(product_12_) );
  ADDFXL U24 ( .A(n84), .B(n88), .CI(n22), .CO(n21), .S(product_11_) );
  ADDFXL U25 ( .A(n89), .B(n91), .CI(n23), .CO(n22), .S(product_10_) );
  ADDFXL U26 ( .A(n93), .B(n92), .CI(n24), .CO(n23), .S(product_9_) );
  ADDFXL U27 ( .A(n94), .B(n97), .CI(n25), .CO(n24), .S(product_8_) );
  ADDFXL U28 ( .A(n98), .B(n99), .CI(n26), .CO(n25), .S(product_7_) );
  ADDFXL U29 ( .A(n100), .B(a_0_), .CI(n27), .CO(n26), .S(product_6_) );
  ADDFXL U30 ( .A(a_1_), .B(n218), .CI(n28), .CO(n27), .S(product_5_) );
  ADDFXL U31 ( .A(a_0_), .B(n219), .CI(n29), .CO(n28), .S(product_4_) );
  ADDHXL U32 ( .A(n220), .B(n30), .CO(n29), .S(product_3_) );
  ADDHXL U33 ( .A(n221), .B(n222), .CO(n30), .S(product_2_) );
  ADDFXL U36 ( .A(n210), .B(n208), .CI(a_15_), .CO(n32), .S(n33) );
  ADDFXL U37 ( .A(n211), .B(a_14_), .CI(n36), .CO(n34), .S(n35) );
  CMPR42X1 U38 ( .A(n212), .B(n210), .C(n209), .D(n207), .ICI(n39), .S(n38), 
        .ICO(n36), .CO(n37) );
  CMPR42X1 U39 ( .A(a_12_), .B(n213), .C(a_14_), .D(n45), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U40 ( .A(n207), .B(n211), .C(n50), .D(n46), .ICI(n47), .S(n44), 
        .ICO(n42), .CO(n43) );
  ADDFXL U41 ( .A(n212), .B(n214), .CI(a_13_), .CO(n45), .S(n46) );
  CMPR42X1 U42 ( .A(n215), .B(a_14_), .C(n51), .D(n55), .ICI(n52), .S(n49), 
        .ICO(n47), .CO(n48) );
  ADDFXL U43 ( .A(n213), .B(a_10_), .CI(a_12_), .CO(n50), .S(n51) );
  CMPR42X1 U44 ( .A(n216), .B(a_13_), .C(n56), .D(n60), .ICI(n57), .S(n54), 
        .ICO(n52), .CO(n53) );
  ADDFXL U45 ( .A(n214), .B(a_9_), .CI(a_11_), .CO(n55), .S(n56) );
  CMPR42X1 U46 ( .A(a_15_), .B(a_12_), .C(n61), .D(n65), .ICI(n62), .S(n59), 
        .ICO(n57), .CO(n58) );
  ADDFXL U47 ( .A(n217), .B(a_8_), .CI(a_10_), .CO(n60), .S(n61) );
  CMPR42X1 U48 ( .A(n208), .B(n215), .C(n70), .D(n66), .ICI(n67), .S(n64), 
        .ICO(n62), .CO(n63) );
  ADDFXL U49 ( .A(a_11_), .B(n218), .CI(a_9_), .CO(n65), .S(n66) );
  CMPR42X1 U50 ( .A(n209), .B(n216), .C(n75), .D(n71), .ICI(n72), .S(n69), 
        .ICO(n67), .CO(n68) );
  ADDFXL U51 ( .A(a_10_), .B(n219), .CI(a_8_), .CO(n70), .S(n71) );
  CMPR42X1 U52 ( .A(n210), .B(n217), .C(n77), .D(n80), .ICI(n76), .S(n74), 
        .ICO(n72), .CO(n73) );
  ADDFXL U53 ( .A(a_9_), .B(n220), .CI(a_7_), .CO(n75), .S(n76) );
  CMPR42X1 U54 ( .A(n211), .B(n218), .C(n85), .D(n82), .ICI(n81), .S(n79), 
        .ICO(n77), .CO(n78) );
  ADDFXL U55 ( .A(a_8_), .B(n221), .CI(a_6_), .CO(n80), .S(n81) );
  CMPR42X1 U56 ( .A(n222), .B(a_5_), .C(a_7_), .D(n87), .ICI(n86), .S(n84), 
        .ICO(n82), .CO(n83) );
  CMPR42X1 U59 ( .A(n213), .B(n220), .C(a_4_), .D(a_6_), .ICI(n90), .S(n89), 
        .ICO(n87), .CO(n88) );
  CMPR42X1 U60 ( .A(n214), .B(n221), .C(a_3_), .D(a_5_), .ICI(n95), .S(n92), 
        .ICO(n90), .CO(n91) );
  ADDFXL U61 ( .A(a_2_), .B(a_4_), .CI(n96), .CO(n93), .S(n94) );
  ADDFXL U64 ( .A(a_1_), .B(n216), .CI(a_3_), .CO(n97), .S(n98) );
  ADDHXL U65 ( .A(n217), .B(a_2_), .CO(n99), .S(n100) );
  CLKINVX1 U87 ( .A(product_28_), .Y(n201) );
  CLKINVX1 U88 ( .A(n201), .Y(product_27_) );
  CLKINVX1 U89 ( .A(n201), .Y(product_29_) );
  CLKINVX1 U90 ( .A(n201), .Y(product_30_) );
  CLKINVX1 U91 ( .A(n201), .Y(product_31_) );
  CLKINVX1 U92 ( .A(a_0_), .Y(n222) );
  CLKINVX1 U93 ( .A(a_2_), .Y(n220) );
  CLKINVX1 U94 ( .A(a_1_), .Y(n221) );
  CLKINVX1 U95 ( .A(a_3_), .Y(n219) );
  CLKINVX1 U96 ( .A(a_7_), .Y(n215) );
  CLKINVX1 U97 ( .A(a_6_), .Y(n216) );
  CLKINVX1 U98 ( .A(a_8_), .Y(n214) );
  CLKINVX1 U99 ( .A(a_5_), .Y(n217) );
  CLKINVX1 U100 ( .A(a_4_), .Y(n218) );
  CLKINVX1 U101 ( .A(a_12_), .Y(n210) );
  CLKINVX1 U102 ( .A(a_10_), .Y(n212) );
  CLKINVX1 U103 ( .A(a_9_), .Y(n213) );
  CLKINVX1 U104 ( .A(a_11_), .Y(n211) );
  CLKINVX1 U105 ( .A(a_14_), .Y(n208) );
  CLKINVX1 U106 ( .A(a_13_), .Y(n209) );
  CLKINVX1 U107 ( .A(a_15_), .Y(n207) );
  CLKBUFX3 U108 ( .A(a_0_), .Y(product_1_) );
  CLKINVX1 U109 ( .A(n6), .Y(product_28_) );
  XOR2X1 U110 ( .A(n215), .B(a_0_), .Y(n96) );
  NAND2X1 U111 ( .A(a_7_), .B(a_0_), .Y(n95) );
  XOR2X1 U112 ( .A(n212), .B(a_3_), .Y(n86) );
  NAND2X1 U113 ( .A(a_10_), .B(a_3_), .Y(n85) );
endmodule


module FIR_FILTER2_DW_mult_uns_4 ( a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_ );
  input a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_,
         a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n172, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195;

  ADDFXL U12 ( .A(a_16_), .B(n182), .CI(n9), .CO(n8), .S(product_24_) );
  ADDFXL U13 ( .A(n29), .B(a_14_), .CI(n10), .CO(n9), .S(product_23_) );
  ADDFXL U14 ( .A(n30), .B(n31), .CI(n11), .CO(n10), .S(product_22_) );
  ADDFXL U15 ( .A(n33), .B(n32), .CI(n12), .CO(n11), .S(product_21_) );
  ADDFXL U16 ( .A(n34), .B(n36), .CI(n13), .CO(n12), .S(product_20_) );
  ADDFXL U17 ( .A(n37), .B(n39), .CI(n14), .CO(n13), .S(product_19_) );
  ADDFXL U18 ( .A(n40), .B(n42), .CI(n15), .CO(n14), .S(product_18_) );
  ADDFXL U19 ( .A(n45), .B(n43), .CI(n16), .CO(n15), .S(product_17_) );
  ADDFXL U20 ( .A(n46), .B(n48), .CI(n17), .CO(n16), .S(product_16_) );
  ADDFXL U21 ( .A(n49), .B(n51), .CI(n18), .CO(n17), .S(product_15_) );
  ADDFXL U22 ( .A(n52), .B(n54), .CI(n19), .CO(n18), .S(product_14_) );
  ADDFXL U23 ( .A(n55), .B(n57), .CI(n20), .CO(n19), .S(product_13_) );
  ADDFXL U24 ( .A(n58), .B(n60), .CI(n21), .CO(n20), .S(product_12_) );
  ADDFXL U25 ( .A(n61), .B(n63), .CI(n22), .CO(n21), .S(product_11_) );
  ADDFXL U26 ( .A(n65), .B(n64), .CI(n23), .CO(n22), .S(product_10_) );
  ADDFXL U27 ( .A(n66), .B(n69), .CI(n24), .CO(n23), .S(product_9_) );
  ADDFXL U28 ( .A(n70), .B(n71), .CI(n25), .CO(n24), .S(product_8_) );
  ADDFXL U29 ( .A(n72), .B(a_5_), .CI(n26), .CO(n25), .S(product_7_) );
  ADDFXL U30 ( .A(a_4_), .B(n194), .CI(n27), .CO(n26), .S(product_6_) );
  ADDFXL U31 ( .A(a_3_), .B(n195), .CI(n28), .CO(n27), .S(product_5_) );
  ADDFXL U34 ( .A(n183), .B(n182), .CI(a_16_), .CO(n29), .S(n30) );
  ADDFXL U35 ( .A(n184), .B(a_14_), .CI(n183), .CO(n31), .S(n32) );
  ADDFXL U36 ( .A(n185), .B(a_13_), .CI(n35), .CO(n33), .S(n34) );
  CMPR42X1 U37 ( .A(n182), .B(n186), .C(n184), .D(a_16_), .ICI(n38), .S(n37), 
        .ICO(n35), .CO(n36) );
  CMPR42X1 U38 ( .A(a_14_), .B(n185), .C(n187), .D(n181), .ICI(n41), .S(n40), 
        .ICO(n38), .CO(n39) );
  CMPR42X1 U39 ( .A(a_15_), .B(n183), .C(n186), .D(n188), .ICI(n44), .S(n43), 
        .ICO(n41), .CO(n42) );
  CMPR42X1 U40 ( .A(n189), .B(n187), .C(n184), .D(a_14_), .ICI(n47), .S(n46), 
        .ICO(n44), .CO(n45) );
  CMPR42X1 U41 ( .A(n190), .B(n188), .C(n185), .D(a_13_), .ICI(n50), .S(n49), 
        .ICO(n47), .CO(n48) );
  CMPR42X1 U42 ( .A(n191), .B(n189), .C(n186), .D(a_12_), .ICI(n53), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U43 ( .A(n192), .B(n190), .C(n187), .D(a_11_), .ICI(n56), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U44 ( .A(n193), .B(n191), .C(n188), .D(a_10_), .ICI(n59), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U45 ( .A(n194), .B(n192), .C(n189), .D(a_9_), .ICI(n62), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U46 ( .A(n195), .B(n193), .C(n190), .D(a_8_), .ICI(n67), .S(n64), 
        .ICO(n62), .CO(n63) );
  ADDFXL U47 ( .A(a_7_), .B(n191), .CI(n68), .CO(n65), .S(n66) );
  ADDFXL U50 ( .A(n192), .B(n195), .CI(a_6_), .CO(n69), .S(n70) );
  CLKINVX1 U77 ( .A(product_28_), .Y(n172) );
  CLKINVX1 U78 ( .A(n172), .Y(product_25_) );
  CLKINVX1 U79 ( .A(n172), .Y(product_26_) );
  CLKINVX1 U80 ( .A(n172), .Y(product_27_) );
  CLKINVX1 U81 ( .A(n172), .Y(product_29_) );
  CLKINVX1 U82 ( .A(n172), .Y(product_30_) );
  CLKINVX1 U83 ( .A(n172), .Y(product_31_) );
  CLKINVX1 U84 ( .A(a_2_), .Y(n194) );
  CLKINVX1 U85 ( .A(a_1_), .Y(n195) );
  CLKINVX1 U86 ( .A(a_6_), .Y(n190) );
  CLKINVX1 U87 ( .A(a_3_), .Y(n193) );
  CLKINVX1 U88 ( .A(a_5_), .Y(n191) );
  CLKINVX1 U89 ( .A(a_4_), .Y(n192) );
  CLKINVX1 U90 ( .A(a_7_), .Y(n189) );
  CLKINVX1 U91 ( .A(a_9_), .Y(n187) );
  CLKINVX1 U92 ( .A(a_8_), .Y(n188) );
  CLKINVX1 U93 ( .A(a_10_), .Y(n186) );
  CLKINVX1 U94 ( .A(a_13_), .Y(n183) );
  CLKINVX1 U95 ( .A(a_11_), .Y(n185) );
  CLKINVX1 U96 ( .A(a_12_), .Y(n184) );
  CLKINVX1 U97 ( .A(a_15_), .Y(n181) );
  CLKINVX1 U98 ( .A(a_14_), .Y(n182) );
  CLKBUFX3 U99 ( .A(a_1_), .Y(product_3_) );
  CLKBUFX3 U100 ( .A(a_0_), .Y(product_2_) );
  XOR2X1 U101 ( .A(a_2_), .B(a_0_), .Y(product_4_) );
  CLKINVX1 U102 ( .A(n8), .Y(product_28_) );
  XOR2X1 U103 ( .A(n193), .B(a_0_), .Y(n72) );
  NAND2X1 U104 ( .A(a_0_), .B(a_3_), .Y(n71) );
  XOR2X1 U105 ( .A(n194), .B(a_0_), .Y(n68) );
  NAND2X1 U106 ( .A(a_0_), .B(a_2_), .Y(n67) );
  NAND2X1 U107 ( .A(a_0_), .B(n194), .Y(n28) );
endmodule


module FIR_FILTER2_DW_mult_uns_3 ( a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_16_, a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_,
         a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114;

  ADDFXL U12 ( .A(a_14_), .B(a_15_), .CI(n9), .CO(product_26_), .S(product_25_) );
  ADDFXL U13 ( .A(n31), .B(a_13_), .CI(n10), .CO(n9), .S(product_24_) );
  ADDFXL U14 ( .A(n32), .B(n34), .CI(n11), .CO(n10), .S(product_23_) );
  ADDFXL U15 ( .A(n35), .B(n37), .CI(n12), .CO(n11), .S(product_22_) );
  ADDFXL U16 ( .A(n38), .B(n40), .CI(n13), .CO(n12), .S(product_21_) );
  ADDFXL U17 ( .A(n43), .B(n41), .CI(n14), .CO(n13), .S(product_20_) );
  ADDFXL U18 ( .A(n44), .B(n46), .CI(n15), .CO(n14), .S(product_19_) );
  ADDFXL U19 ( .A(n47), .B(n51), .CI(n16), .CO(n15), .S(product_18_) );
  ADDFXL U20 ( .A(n52), .B(n57), .CI(n17), .CO(n16), .S(product_17_) );
  ADDFXL U21 ( .A(n58), .B(n63), .CI(n18), .CO(n17), .S(product_16_) );
  ADDFXL U22 ( .A(n64), .B(n69), .CI(n19), .CO(n18), .S(product_15_) );
  ADDFXL U23 ( .A(n70), .B(n75), .CI(n20), .CO(n19), .S(product_14_) );
  ADDFXL U24 ( .A(n76), .B(n81), .CI(n21), .CO(n20), .S(product_13_) );
  ADDFXL U25 ( .A(n82), .B(n87), .CI(n22), .CO(n21), .S(product_12_) );
  ADDFXL U26 ( .A(n88), .B(n94), .CI(n23), .CO(n22), .S(product_11_) );
  ADDFXL U27 ( .A(n95), .B(n99), .CI(n24), .CO(n23), .S(product_10_) );
  ADDFXL U28 ( .A(n103), .B(n100), .CI(n25), .CO(n24), .S(product_9_) );
  ADDFXL U29 ( .A(n104), .B(n107), .CI(n26), .CO(n25), .S(product_8_) );
  ADDFXL U30 ( .A(n108), .B(n109), .CI(n27), .CO(n26), .S(product_7_) );
  ADDFXL U31 ( .A(n110), .B(n111), .CI(n28), .CO(n27), .S(product_6_) );
  ADDFXL U32 ( .A(n112), .B(n113), .CI(n29), .CO(n28), .S(product_5_) );
  ADDFXL U33 ( .A(n91), .B(a_0_), .CI(n114), .CO(n29), .S(product_4_) );
  ADDFXL U35 ( .A(a_12_), .B(a_14_), .CI(n33), .CO(n31), .S(n32) );
  CMPR42X1 U36 ( .A(a_15_), .B(a_14_), .C(a_11_), .D(a_13_), .ICI(n36), .S(n35), .ICO(n33), .CO(n34) );
  CMPR42X1 U37 ( .A(a_15_), .B(a_13_), .C(a_10_), .D(a_12_), .ICI(n39), .S(n38), .ICO(n36), .CO(n37) );
  CMPR42X1 U38 ( .A(a_15_), .B(a_12_), .C(a_9_), .D(a_11_), .ICI(n42), .S(n41), 
        .ICO(n39), .CO(n40) );
  CMPR42X1 U39 ( .A(a_11_), .B(a_8_), .C(a_10_), .D(n48), .ICI(n45), .S(n44), 
        .ICO(n42), .CO(n43) );
  CMPR42X1 U40 ( .A(a_9_), .B(n53), .C(n54), .D(n49), .ICI(n50), .S(n47), 
        .ICO(n45), .CO(n46) );
  ADDFXL U41 ( .A(a_10_), .B(a_14_), .CI(a_7_), .CO(n48), .S(n49) );
  CMPR42X1 U42 ( .A(a_13_), .B(n59), .C(n60), .D(n55), .ICI(n56), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U43 ( .A(a_15_), .B(a_8_), .C(a_6_), .D(a_14_), .ICI(a_9_), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U44 ( .A(a_12_), .B(n65), .C(n61), .D(n66), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U45 ( .A(a_15_), .B(a_7_), .C(a_5_), .D(a_13_), .ICI(a_8_), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U46 ( .A(a_12_), .B(a_11_), .C(n72), .D(n67), .ICI(n68), .S(n64), 
        .ICO(n62), .CO(n63) );
  CMPR42X1 U47 ( .A(a_6_), .B(a_4_), .C(a_7_), .D(a_14_), .ICI(n71), .S(n67), 
        .ICO(n65), .CO(n66) );
  CMPR42X1 U48 ( .A(a_11_), .B(a_10_), .C(n78), .D(n73), .ICI(n74), .S(n70), 
        .ICO(n68), .CO(n69) );
  CMPR42X1 U49 ( .A(a_5_), .B(a_3_), .C(a_6_), .D(a_13_), .ICI(n77), .S(n73), 
        .ICO(n71), .CO(n72) );
  CMPR42X1 U50 ( .A(a_10_), .B(a_9_), .C(n84), .D(n79), .ICI(n80), .S(n76), 
        .ICO(n74), .CO(n75) );
  CMPR42X1 U51 ( .A(a_4_), .B(a_2_), .C(a_5_), .D(a_12_), .ICI(n83), .S(n79), 
        .ICO(n77), .CO(n78) );
  CMPR42X1 U52 ( .A(a_11_), .B(a_9_), .C(n89), .D(n85), .ICI(n86), .S(n82), 
        .ICO(n80), .CO(n81) );
  CMPR42X1 U53 ( .A(a_3_), .B(a_1_), .C(a_4_), .D(a_8_), .ICI(n91), .S(n85), 
        .ICO(n83), .CO(n84) );
  CMPR42X1 U54 ( .A(a_10_), .B(product_3_), .C(n93), .D(n96), .ICI(n90), .S(
        n88), .ICO(n86), .CO(n87) );
  ADDFXL U55 ( .A(a_3_), .B(a_7_), .CI(a_8_), .CO(n89), .S(n90) );
  ADDHXL U56 ( .A(a_2_), .B(a_0_), .CO(n91), .S(product_3_) );
  CMPR42X1 U57 ( .A(a_9_), .B(a_7_), .C(n101), .D(n98), .ICI(n97), .S(n95), 
        .ICO(n93), .CO(n94) );
  ADDFXL U58 ( .A(a_1_), .B(a_2_), .CI(a_6_), .CO(n96), .S(n97) );
  CMPR42X1 U59 ( .A(a_8_), .B(a_5_), .C(a_6_), .D(n105), .ICI(n102), .S(n100), 
        .ICO(n98), .CO(n99) );
  ADDHXL U60 ( .A(a_1_), .B(a_0_), .CO(n101), .S(n102) );
  ADDFXL U61 ( .A(a_5_), .B(a_7_), .CI(n106), .CO(n103), .S(n104) );
  ADDHXL U62 ( .A(a_4_), .B(a_0_), .CO(n105), .S(n106) );
  ADDFXL U63 ( .A(a_3_), .B(a_6_), .CI(a_4_), .CO(n107), .S(n108) );
  ADDFXL U64 ( .A(a_2_), .B(a_5_), .CI(a_3_), .CO(n109), .S(n110) );
  ADDFXL U65 ( .A(a_1_), .B(a_4_), .CI(a_2_), .CO(n111), .S(n112) );
  ADDHXL U66 ( .A(a_3_), .B(a_1_), .CO(n113), .S(n114) );
  CLKBUFX3 U87 ( .A(a_16_), .Y(product_27_) );
  CLKBUFX3 U88 ( .A(a_16_), .Y(product_28_) );
  CLKBUFX3 U89 ( .A(a_16_), .Y(product_29_) );
  CLKBUFX3 U90 ( .A(a_16_), .Y(product_30_) );
  CLKBUFX3 U91 ( .A(a_16_), .Y(product_31_) );
  CLKBUFX3 U92 ( .A(a_1_), .Y(product_2_) );
  CLKBUFX3 U93 ( .A(a_0_), .Y(product_1_) );
endmodule


module FIR_FILTER2_DW_mult_uns_2 ( a_16_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_ );
  input a_16_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211;

  ADDFXL U5 ( .A(a_14_), .B(n196), .CI(n4), .CO(n3), .S(product_28_) );
  ADDFXL U6 ( .A(n197), .B(a_13_), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U7 ( .A(n198), .B(a_12_), .CI(n6), .CO(n5), .S(product_26_) );
  ADDFXL U8 ( .A(n36), .B(n199), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U9 ( .A(n37), .B(n38), .CI(n8), .CO(n7), .S(product_24_) );
  ADDFXL U10 ( .A(n40), .B(n39), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U11 ( .A(n41), .B(n43), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U12 ( .A(n46), .B(n44), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U13 ( .A(n47), .B(n49), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U14 ( .A(n50), .B(n54), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U15 ( .A(n55), .B(n59), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U16 ( .A(n60), .B(n64), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U17 ( .A(n65), .B(n69), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U18 ( .A(n70), .B(n74), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U19 ( .A(n75), .B(n79), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U20 ( .A(n80), .B(n84), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U21 ( .A(n85), .B(n89), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U22 ( .A(n90), .B(n94), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U23 ( .A(n95), .B(n99), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U24 ( .A(n101), .B(n100), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U25 ( .A(n102), .B(n105), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U26 ( .A(n106), .B(n109), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U27 ( .A(n110), .B(n111), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFXL U28 ( .A(n112), .B(n209), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFXL U29 ( .A(n211), .B(a_2_), .CI(n28), .CO(n27), .S(product_4_) );
  ADDHXL U30 ( .A(n210), .B(n211), .CO(n28), .S(product_3_) );
  ADDFXL U36 ( .A(a_11_), .B(n197), .CI(a_16_), .CO(n36), .S(n37) );
  ADDFXL U37 ( .A(n198), .B(a_14_), .CI(a_10_), .CO(n38), .S(n39) );
  ADDFXL U38 ( .A(a_9_), .B(a_13_), .CI(n42), .CO(n40), .S(n41) );
  CMPR42X1 U39 ( .A(n197), .B(n199), .C(a_8_), .D(a_16_), .ICI(n45), .S(n44), 
        .ICO(n42), .CO(n43) );
  CMPR42X1 U40 ( .A(a_14_), .B(n200), .C(a_7_), .D(n51), .ICI(n48), .S(n47), 
        .ICO(n45), .CO(n46) );
  CMPR42X1 U41 ( .A(n198), .B(n201), .C(n56), .D(n52), .ICI(n53), .S(n50), 
        .ICO(n48), .CO(n49) );
  ADDFXL U42 ( .A(a_6_), .B(n197), .CI(a_16_), .CO(n51), .S(n52) );
  CMPR42X1 U43 ( .A(n199), .B(n202), .C(n61), .D(n57), .ICI(n58), .S(n55), 
        .ICO(n53), .CO(n54) );
  ADDFXL U44 ( .A(n198), .B(a_14_), .CI(a_5_), .CO(n56), .S(n57) );
  CMPR42X1 U45 ( .A(n203), .B(a_16_), .C(n62), .D(n66), .ICI(n63), .S(n60), 
        .ICO(n58), .CO(n59) );
  ADDFXL U46 ( .A(n200), .B(a_13_), .CI(a_4_), .CO(n61), .S(n62) );
  CMPR42X1 U47 ( .A(n199), .B(n201), .C(n71), .D(n67), .ICI(n68), .S(n65), 
        .ICO(n63), .CO(n64) );
  ADDFXL U48 ( .A(n204), .B(n197), .CI(a_3_), .CO(n66), .S(n67) );
  CMPR42X1 U49 ( .A(n200), .B(n202), .C(n76), .D(n72), .ICI(n73), .S(n70), 
        .ICO(n68), .CO(n69) );
  ADDFXL U50 ( .A(n205), .B(n198), .CI(a_2_), .CO(n71), .S(n72) );
  CMPR42X1 U51 ( .A(n201), .B(n203), .C(n78), .D(n81), .ICI(n77), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U52 ( .A(n206), .B(n199), .CI(a_1_), .CO(n76), .S(n77) );
  CMPR42X1 U53 ( .A(n202), .B(n204), .C(n86), .D(n83), .ICI(n82), .S(n80), 
        .ICO(n78), .CO(n79) );
  ADDFXL U54 ( .A(n207), .B(n200), .CI(a_0_), .CO(n81), .S(n82) );
  CMPR42X1 U55 ( .A(n201), .B(n203), .C(n91), .D(n87), .ICI(n88), .S(n85), 
        .ICO(n83), .CO(n84) );
  ADDHXL U56 ( .A(n205), .B(n208), .CO(n86), .S(n87) );
  CMPR42X1 U57 ( .A(n202), .B(n204), .C(n96), .D(n93), .ICI(n92), .S(n90), 
        .ICO(n88), .CO(n89) );
  ADDHXL U58 ( .A(n206), .B(n209), .CO(n91), .S(n92) );
  CMPR42X1 U59 ( .A(n203), .B(n207), .C(n205), .D(n98), .ICI(n97), .S(n95), 
        .ICO(n93), .CO(n94) );
  ADDHXL U60 ( .A(n210), .B(n204), .CO(n96), .S(n97) );
  CMPR42X1 U61 ( .A(a_7_), .B(n206), .C(n211), .D(n208), .ICI(n103), .S(n100), 
        .ICO(n98), .CO(n99) );
  ADDFXL U62 ( .A(n107), .B(n207), .CI(n104), .CO(n101), .S(n102) );
  ADDHXL U63 ( .A(n205), .B(n209), .CO(n103), .S(n104) );
  ADDFXL U64 ( .A(n208), .B(n206), .CI(n108), .CO(n105), .S(n106) );
  ADDHXL U65 ( .A(n210), .B(n207), .CO(n107), .S(n108) );
  ADDFXL U66 ( .A(n211), .B(a_4_), .CI(n209), .CO(n109), .S(n110) );
  ADDHXL U67 ( .A(n208), .B(n210), .CO(n111), .S(n112) );
  CLKBUFX3 U91 ( .A(product_29_), .Y(product_30_) );
  CLKBUFX3 U92 ( .A(product_29_), .Y(product_31_) );
  CLKINVX1 U93 ( .A(a_16_), .Y(n196) );
  CLKINVX1 U94 ( .A(a_4_), .Y(n207) );
  CLKINVX1 U95 ( .A(a_0_), .Y(n211) );
  CLKINVX1 U96 ( .A(a_2_), .Y(n209) );
  CLKINVX1 U97 ( .A(a_5_), .Y(n206) );
  CLKINVX1 U98 ( .A(a_3_), .Y(n208) );
  CLKINVX1 U99 ( .A(a_6_), .Y(n205) );
  CLKINVX1 U100 ( .A(a_1_), .Y(n210) );
  CLKINVX1 U101 ( .A(a_8_), .Y(n203) );
  CLKINVX1 U102 ( .A(a_9_), .Y(n202) );
  CLKINVX1 U103 ( .A(a_7_), .Y(n204) );
  CLKINVX1 U104 ( .A(a_12_), .Y(n199) );
  CLKINVX1 U105 ( .A(a_14_), .Y(n197) );
  CLKINVX1 U106 ( .A(a_10_), .Y(n201) );
  CLKINVX1 U107 ( .A(a_13_), .Y(n198) );
  CLKINVX1 U108 ( .A(a_11_), .Y(n200) );
  CLKBUFX3 U109 ( .A(a_0_), .Y(product_2_) );
  CLKINVX1 U110 ( .A(n3), .Y(product_29_) );
endmodule


module FIR_FILTER2_DW_mult_uns_1 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_
 );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n34, n35,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201;

  ADDFXL U5 ( .A(a_14_), .B(n186), .CI(n4), .CO(n3), .S(product_28_) );
  ADDFXL U6 ( .A(a_13_), .B(n186), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U7 ( .A(n187), .B(a_12_), .CI(n6), .CO(n5), .S(product_26_) );
  ADDFXL U8 ( .A(n188), .B(a_11_), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U9 ( .A(n34), .B(n189), .CI(n8), .CO(n7), .S(product_24_) );
  ADDFXL U10 ( .A(n35), .B(n38), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U11 ( .A(n41), .B(n39), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U12 ( .A(n42), .B(n44), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U13 ( .A(n45), .B(n49), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U14 ( .A(n50), .B(n54), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U15 ( .A(n55), .B(n59), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U16 ( .A(n60), .B(n64), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U17 ( .A(n65), .B(n69), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U18 ( .A(n70), .B(n74), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U19 ( .A(n75), .B(n79), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U20 ( .A(n83), .B(n80), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U21 ( .A(n84), .B(n87), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U22 ( .A(n88), .B(n89), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U23 ( .A(n90), .B(n91), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U24 ( .A(n92), .B(n93), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U25 ( .A(n94), .B(n95), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U26 ( .A(n96), .B(a_2_), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U27 ( .A(a_1_), .B(n196), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFXL U28 ( .A(a_0_), .B(n197), .CI(n27), .CO(n26), .S(product_5_) );
  ADDHXL U29 ( .A(n198), .B(n28), .CO(n27), .S(product_4_) );
  ADDHXL U30 ( .A(n199), .B(n29), .CO(n28), .S(product_3_) );
  ADDHXL U31 ( .A(n200), .B(n201), .CO(n29), .S(product_2_) );
  ADDFXL U36 ( .A(n190), .B(a_10_), .CI(n37), .CO(n34), .S(n35) );
  CMPR42X1 U38 ( .A(n187), .B(a_9_), .C(a_10_), .D(a_15_), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U39 ( .A(a_14_), .B(a_9_), .C(a_8_), .D(n46), .ICI(n43), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U40 ( .A(n186), .B(n188), .C(n51), .D(n47), .ICI(n48), .S(n45), 
        .ICO(n43), .CO(n44) );
  ADDFXL U41 ( .A(a_8_), .B(n189), .CI(a_7_), .CO(n46), .S(n47) );
  CMPR42X1 U42 ( .A(a_14_), .B(a_7_), .C(n56), .D(n52), .ICI(n53), .S(n50), 
        .ICO(n48), .CO(n49) );
  ADDFXL U43 ( .A(n190), .B(a_12_), .CI(a_6_), .CO(n51), .S(n52) );
  CMPR42X1 U44 ( .A(a_13_), .B(a_6_), .C(n61), .D(n57), .ICI(n58), .S(n55), 
        .ICO(n53), .CO(n54) );
  ADDFXL U45 ( .A(n191), .B(a_11_), .CI(a_5_), .CO(n56), .S(n57) );
  CMPR42X1 U46 ( .A(a_12_), .B(a_5_), .C(n62), .D(n66), .ICI(n63), .S(n60), 
        .ICO(n58), .CO(n59) );
  ADDFXL U47 ( .A(n192), .B(a_10_), .CI(a_4_), .CO(n61), .S(n62) );
  CMPR42X1 U48 ( .A(a_15_), .B(a_11_), .C(n67), .D(n71), .ICI(n68), .S(n65), 
        .ICO(n63), .CO(n64) );
  ADDFXL U49 ( .A(a_4_), .B(a_9_), .CI(a_3_), .CO(n66), .S(n67) );
  CMPR42X1 U50 ( .A(n193), .B(a_10_), .C(n73), .D(n76), .ICI(n72), .S(n70), 
        .ICO(n68), .CO(n69) );
  ADDFXL U51 ( .A(a_2_), .B(n187), .CI(a_3_), .CO(n71), .S(n72) );
  CMPR42X1 U52 ( .A(n194), .B(a_9_), .C(n81), .D(n78), .ICI(n77), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U53 ( .A(a_1_), .B(n188), .CI(a_2_), .CO(n76), .S(n77) );
  CMPR42X1 U54 ( .A(n195), .B(a_1_), .C(a_8_), .D(n85), .ICI(n82), .S(n80), 
        .ICO(n78), .CO(n79) );
  ADDHXL U55 ( .A(n189), .B(a_0_), .CO(n81), .S(n82) );
  ADDFXL U56 ( .A(a_7_), .B(n196), .CI(n86), .CO(n83), .S(n84) );
  ADDHXL U57 ( .A(n190), .B(a_0_), .CO(n85), .S(n86) );
  ADDFXL U58 ( .A(n197), .B(n191), .CI(a_6_), .CO(n87), .S(n88) );
  ADDFXL U59 ( .A(n198), .B(n192), .CI(a_5_), .CO(n89), .S(n90) );
  ADDFXL U60 ( .A(n199), .B(n193), .CI(a_4_), .CO(n91), .S(n92) );
  ADDFXL U61 ( .A(n200), .B(n194), .CI(a_3_), .CO(n93), .S(n94) );
  CLKBUFX3 U89 ( .A(product_29_), .Y(product_30_) );
  CLKBUFX3 U90 ( .A(product_29_), .Y(product_31_) );
  CLKINVX1 U91 ( .A(a_0_), .Y(n201) );
  CLKINVX1 U92 ( .A(a_7_), .Y(n194) );
  CLKINVX1 U93 ( .A(a_5_), .Y(n196) );
  CLKINVX1 U94 ( .A(a_1_), .Y(n200) );
  CLKINVX1 U95 ( .A(a_3_), .Y(n198) );
  CLKINVX1 U96 ( .A(a_4_), .Y(n197) );
  CLKINVX1 U97 ( .A(a_2_), .Y(n199) );
  CLKINVX1 U98 ( .A(a_6_), .Y(n195) );
  CLKINVX1 U99 ( .A(a_9_), .Y(n192) );
  CLKINVX1 U100 ( .A(a_8_), .Y(n193) );
  CLKINVX1 U101 ( .A(a_10_), .Y(n191) );
  CLKINVX1 U102 ( .A(a_14_), .Y(n187) );
  CLKINVX1 U103 ( .A(a_13_), .Y(n188) );
  CLKINVX1 U104 ( .A(a_12_), .Y(n189) );
  CLKINVX1 U105 ( .A(a_11_), .Y(n190) );
  CLKINVX1 U106 ( .A(a_15_), .Y(n186) );
  CLKBUFX3 U107 ( .A(a_0_), .Y(product_1_) );
  CLKINVX1 U108 ( .A(n3), .Y(product_29_) );
  XOR2X1 U109 ( .A(n195), .B(a_0_), .Y(n96) );
  NAND2X1 U110 ( .A(a_6_), .B(a_0_), .Y(n95) );
endmodule


module FIR_FILTER2_DW_mult_uns_0 ( a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, 
        a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        product_31_, product_30_, product_29_, product_28_, product_27_, 
        product_26_, product_25_, product_24_, product_23_, product_22_, 
        product_21_, product_20_, product_19_, product_18_, product_17_, 
        product_16_, product_15_, product_14_, product_13_, product_12_, 
        product_11_, product_10_, product_9_, product_8_, product_7_, 
        product_6_, product_5_, product_4_, product_3_, product_2_, product_1_, 
        product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259;

  ADDFXL U4 ( .A(a_14_), .B(n245), .CI(n3), .CO(n2), .S(product_29_) );
  ADDFXL U5 ( .A(n246), .B(a_13_), .CI(n4), .CO(n3), .S(product_28_) );
  ADDFXL U6 ( .A(n33), .B(n247), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U7 ( .A(n34), .B(n35), .CI(n6), .CO(n5), .S(product_26_) );
  ADDFXL U8 ( .A(n36), .B(n38), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U9 ( .A(n41), .B(n39), .CI(n8), .CO(n7), .S(product_24_) );
  ADDFXL U10 ( .A(n42), .B(n44), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U11 ( .A(n45), .B(n49), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U12 ( .A(n50), .B(n54), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U13 ( .A(n60), .B(n55), .CI(n12), .CO(n11), .S(product_20_) );
  ADDFXL U14 ( .A(n66), .B(n61), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U15 ( .A(n67), .B(n74), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U16 ( .A(n75), .B(n82), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFXL U17 ( .A(n83), .B(n90), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFXL U18 ( .A(n91), .B(n98), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFXL U19 ( .A(n99), .B(n106), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFXL U20 ( .A(n107), .B(n112), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFXL U21 ( .A(n113), .B(n118), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFXL U22 ( .A(n119), .B(n125), .CI(n21), .CO(n20), .S(product_11_) );
  ADDFXL U23 ( .A(n126), .B(n130), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFXL U24 ( .A(n131), .B(n135), .CI(n23), .CO(n22), .S(product_9_) );
  ADDFXL U25 ( .A(n137), .B(n136), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFXL U26 ( .A(n138), .B(n141), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFXL U27 ( .A(n142), .B(n143), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFXL U28 ( .A(n144), .B(a_0_), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFXL U29 ( .A(a_4_), .B(a_1_), .CI(n28), .CO(n27), .S(product_4_) );
  ADDHXL U30 ( .A(a_0_), .B(a_3_), .CO(n28), .S(product_3_) );
  ADDFXL U35 ( .A(a_12_), .B(n246), .CI(a_15_), .CO(n33), .S(n34) );
  ADDFXL U36 ( .A(a_11_), .B(a_14_), .CI(n37), .CO(n35), .S(n36) );
  CMPR42X1 U37 ( .A(n245), .B(n248), .C(n247), .D(a_10_), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U38 ( .A(a_12_), .B(a_14_), .C(a_9_), .D(n46), .ICI(n43), .S(n42), 
        .ICO(n40), .CO(n41) );
  CMPR42X1 U39 ( .A(n245), .B(n249), .C(n51), .D(n47), .ICI(n48), .S(n45), 
        .ICO(n43), .CO(n44) );
  ADDFXL U40 ( .A(a_13_), .B(n250), .CI(a_8_), .CO(n46), .S(n47) );
  CMPR42X1 U41 ( .A(a_14_), .B(n56), .C(n52), .D(n57), .ICI(n53), .S(n50), 
        .ICO(n48), .CO(n49) );
  ADDFXL U42 ( .A(a_12_), .B(a_10_), .CI(a_7_), .CO(n51), .S(n52) );
  CMPR42X1 U43 ( .A(n245), .B(n251), .C(n63), .D(n58), .ICI(n59), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U44 ( .A(n252), .B(a_6_), .C(a_11_), .D(a_13_), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U45 ( .A(a_5_), .B(n71), .C(n69), .D(n64), .ICI(n65), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U46 ( .A(a_8_), .B(a_10_), .C(a_14_), .D(a_12_), .ICI(n68), .S(n64), 
        .ICO(n62), .CO(n63) );
  CMPR42X1 U47 ( .A(n79), .B(n72), .C(n77), .D(n70), .ICI(n73), .S(n67), .ICO(
        n65), .CO(n66) );
  CMPR42X1 U48 ( .A(n245), .B(n253), .C(a_13_), .D(a_11_), .ICI(n76), .S(n70), 
        .ICO(n68), .CO(n69) );
  ADDFXL U49 ( .A(a_4_), .B(n254), .CI(a_9_), .CO(n71), .S(n72) );
  CMPR42X1 U50 ( .A(n87), .B(n80), .C(n85), .D(n78), .ICI(n81), .S(n75), .ICO(
        n73), .CO(n74) );
  CMPR42X1 U51 ( .A(a_8_), .B(a_12_), .C(a_10_), .D(a_3_), .ICI(n84), .S(n78), 
        .ICO(n76), .CO(n77) );
  ADDFXL U52 ( .A(n255), .B(a_6_), .CI(a_14_), .CO(n79), .S(n80) );
  CMPR42X1 U53 ( .A(n95), .B(n88), .C(n93), .D(n86), .ICI(n89), .S(n83), .ICO(
        n81), .CO(n82) );
  CMPR42X1 U54 ( .A(a_7_), .B(a_11_), .C(a_9_), .D(a_2_), .ICI(n92), .S(n86), 
        .ICO(n84), .CO(n85) );
  ADDFXL U55 ( .A(n245), .B(a_5_), .CI(a_13_), .CO(n87), .S(n88) );
  CMPR42X1 U56 ( .A(n103), .B(n96), .C(n101), .D(n94), .ICI(n97), .S(n91), 
        .ICO(n89), .CO(n90) );
  CMPR42X1 U57 ( .A(a_12_), .B(a_6_), .C(a_10_), .D(a_8_), .ICI(n100), .S(n94), 
        .ICO(n92), .CO(n93) );
  ADDFXL U58 ( .A(n256), .B(a_15_), .CI(a_1_), .CO(n95), .S(n96) );
  CMPR42X1 U59 ( .A(a_9_), .B(n104), .C(n109), .D(n102), .ICI(n105), .S(n99), 
        .ICO(n97), .CO(n98) );
  CMPR42X1 U60 ( .A(a_14_), .B(a_5_), .C(a_11_), .D(a_7_), .ICI(n108), .S(n102), .ICO(n100), .CO(n101) );
  ADDHXL U61 ( .A(n257), .B(a_0_), .CO(n103), .S(n104) );
  CMPR42X1 U62 ( .A(a_10_), .B(a_8_), .C(n115), .D(n110), .ICI(n111), .S(n107), 
        .ICO(n105), .CO(n106) );
  CMPR42X1 U63 ( .A(n258), .B(a_4_), .C(a_6_), .D(a_13_), .ICI(n114), .S(n110), 
        .ICO(n108), .CO(n109) );
  CMPR42X1 U64 ( .A(a_12_), .B(a_9_), .C(n120), .D(n116), .ICI(n117), .S(n113), 
        .ICO(n111), .CO(n112) );
  CMPR42X1 U65 ( .A(n259), .B(a_3_), .C(a_5_), .D(a_7_), .ICI(n122), .S(n116), 
        .ICO(n114), .CO(n115) );
  CMPR42X1 U66 ( .A(a_11_), .B(n123), .C(n124), .D(n127), .ICI(n121), .S(n119), 
        .ICO(n117), .CO(n118) );
  ADDFXL U67 ( .A(a_2_), .B(a_6_), .CI(a_8_), .CO(n120), .S(n121) );
  CMPR42X1 U70 ( .A(a_10_), .B(a_7_), .C(n139), .D(n129), .ICI(n128), .S(n126), 
        .ICO(n124), .CO(n125) );
  ADDFXL U71 ( .A(a_1_), .B(a_3_), .CI(a_5_), .CO(n127), .S(n128) );
  CMPR42X1 U72 ( .A(a_9_), .B(a_4_), .C(a_6_), .D(n134), .ICI(n140), .S(n131), 
        .ICO(n129), .CO(n130) );
  CMPR42X1 U74 ( .A(a_3_), .B(a_1_), .C(a_5_), .D(a_8_), .ICI(n139), .S(n136), 
        .ICO(n134), .CO(n135) );
  ADDFXL U75 ( .A(a_4_), .B(a_7_), .CI(n140), .CO(n137), .S(n138) );
  ADDHXL U76 ( .A(a_2_), .B(a_0_), .CO(n139), .S(n140) );
  ADDFXL U77 ( .A(a_1_), .B(a_6_), .CI(a_3_), .CO(n141), .S(n142) );
  ADDHXL U78 ( .A(a_5_), .B(a_2_), .CO(n143), .S(n144) );
  CLKBUFX3 U114 ( .A(product_31_), .Y(product_30_) );
  CLKINVX1 U115 ( .A(a_1_), .Y(n259) );
  CLKINVX1 U116 ( .A(a_2_), .Y(n258) );
  CLKINVX1 U117 ( .A(a_4_), .Y(n256) );
  CLKINVX1 U118 ( .A(a_3_), .Y(n257) );
  INVX3 U119 ( .A(a_15_), .Y(n245) );
  CLKINVX1 U120 ( .A(a_5_), .Y(n255) );
  CLKINVX1 U121 ( .A(a_6_), .Y(n254) );
  CLKINVX1 U122 ( .A(a_7_), .Y(n253) );
  CLKINVX1 U123 ( .A(a_8_), .Y(n252) );
  CLKINVX1 U124 ( .A(a_9_), .Y(n251) );
  CLKINVX1 U125 ( .A(a_10_), .Y(n250) );
  CLKINVX1 U126 ( .A(a_11_), .Y(n249) );
  CLKINVX1 U127 ( .A(a_12_), .Y(n248) );
  CLKINVX1 U128 ( .A(a_13_), .Y(n247) );
  CLKINVX1 U129 ( .A(a_14_), .Y(n246) );
  CLKBUFX3 U130 ( .A(a_1_), .Y(product_1_) );
  CLKBUFX3 U131 ( .A(a_0_), .Y(product_0_) );
  CLKBUFX3 U132 ( .A(a_2_), .Y(product_2_) );
  CLKINVX1 U133 ( .A(n2), .Y(product_31_) );
  XOR2X1 U134 ( .A(a_4_), .B(a_0_), .Y(n123) );
  NAND2X1 U135 ( .A(a_0_), .B(n256), .Y(n122) );
endmodule


module FIR_FILTER2 ( clk, rst, data_valid, data, fir_valid, fir_d );
  input [15:0] data;
  output [15:0] fir_d;
  input clk, rst, data_valid;
  output fir_valid;
  wire   n149, N7, N12, N13, N14, N15, N16, N17, N20, N21, N22, N23, N24, N54,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n701, n71, n72, N99, N98, N97, N96, N95, N94, N93,
         N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79,
         N78, N77, N76, N75, N74, N73, N720, N710, N702, N690, N680, N670,
         N660, N650, N640, N630, N620, N610, N600, N590, N580, N57, N503, N502,
         N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491,
         N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480,
         N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469,
         N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458,
         N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447,
         N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436,
         N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425,
         N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414,
         N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403,
         N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392,
         N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381,
         N380, N379, N378, N377, N375, N374, N373, N372, N371, N370, N369,
         N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358,
         N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347,
         N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336,
         N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325,
         N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314,
         N313, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302,
         N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291,
         N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280,
         N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269,
         N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258,
         N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247,
         N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236,
         N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225,
         N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214,
         N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203,
         N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192,
         N191, N190, N189, N188, N187, N186, N185, N183, N182, N181, N180,
         N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169,
         N168, N167, N166, N165, N164, N163, N162, N161, N1600, N159, N158,
         N157, N156, N155, N154, N153, N152, N151, N1500, N1490, N148, N147,
         N146, N145, N144, N143, N142, N141, N1401, N139, N138, N137, N136,
         N135, N134, N133, N132, N131, N1301, N129, N128, N127, N126, N125,
         N124, N123, N122, N121, N1201, N119, N118, N117, N116, N115, N114,
         N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103,
         N102, N101, N100, mult_120_n29, mult_120_n28, mult_120_n27,
         mult_120_n26, mult_120_n25, mult_120_n24, mult_120_n23, mult_120_n22,
         mult_120_n21, mult_120_n20, mult_120_n19, mult_120_n18, mult_120_n17,
         mult_120_n16, mult_120_n15, mult_120_n14, n18, n19, n2010, n2110,
         n2210, n2310, n2410, n25, n26, n27, n28, n29, n30, n31, n32, n33, n50,
         n53, n540, n55, n56, n570, n730, n740, n750, n760, n770, n780, n790,
         n800, n810, n820, n830, n840, n850, n860, n870, n880, n890, n900,
         n910, n920, n930, n940, n950, n960, n970, n980, n990, n1000, n1010,
         n1020, n1030;
  wire   [5:0] cnt_data;
  wire   [511:0] fir_data;
  wire   [255:0] add_fir;
  wire   [252:0] temp_add_fir;
  wire   [487:0] mul_add_fir;
  wire   [511:0] temp_mul_add_fir;
  wire   [31:16] comb_fir_o;
  wire   [15:0] revise_o;
  wire   [5:2] add_55_carry;

  DFFRX4 fir_d_reg_14_ ( .D(revise_o[14]), .CK(clk), .RN(n1030), .QN(n32) );
  DFFRX4 fir_d_reg_13_ ( .D(revise_o[13]), .CK(clk), .RN(n1030), .QN(n31) );
  DFFRX4 fir_d_reg_12_ ( .D(revise_o[12]), .CK(clk), .RN(n1030), .QN(n30) );
  DFFRX4 fir_d_reg_11_ ( .D(revise_o[11]), .CK(clk), .RN(n1030), .QN(n29) );
  DFFRX4 fir_d_reg_10_ ( .D(revise_o[10]), .CK(clk), .RN(n1030), .QN(n28) );
  DFFRX4 fir_d_reg_9_ ( .D(revise_o[9]), .CK(clk), .RN(n1030), .QN(n27) );
  DFFRX4 fir_d_reg_8_ ( .D(revise_o[8]), .CK(clk), .RN(n1030), .QN(n26) );
  DFFRX4 fir_d_reg_7_ ( .D(revise_o[7]), .CK(clk), .RN(n1030), .QN(n2210) );
  DFFRX4 fir_d_reg_6_ ( .D(revise_o[6]), .CK(clk), .RN(n1030), .QN(n2310) );
  DFFRX4 fir_d_reg_5_ ( .D(revise_o[5]), .CK(clk), .RN(n1030), .QN(n25) );
  DFFRX4 fir_d_reg_4_ ( .D(revise_o[4]), .CK(clk), .RN(n1030), .QN(n2410) );
  DFFRX4 fir_d_reg_3_ ( .D(revise_o[3]), .CK(clk), .RN(n1030), .QN(n2110) );
  DFFRX4 fir_d_reg_2_ ( .D(revise_o[2]), .CK(clk), .RN(n1030), .QN(n2010) );
  DFFRX4 fir_d_reg_1_ ( .D(revise_o[1]), .CK(clk), .RN(n1030), .QN(n19) );
  DFFRX4 fir_d_reg_0_ ( .D(revise_o[0]), .CK(clk), .RN(n1030), .QN(n18) );
  FIR_FILTER2_DW01_add_0 add_111 ( .A(fir_data[271:256]), .B(fir_data[255:240]), .SUM(add_fir[15:0]) );
  FIR_FILTER2_DW01_add_1 add_110 ( .A(fir_data[287:272]), .B(fir_data[239:224]), .SUM(add_fir[31:16]) );
  FIR_FILTER2_DW01_add_2 add_109 ( .A(fir_data[303:288]), .B(fir_data[223:208]), .SUM(add_fir[47:32]) );
  FIR_FILTER2_DW01_add_3 add_108 ( .A(fir_data[319:304]), .B(fir_data[207:192]), .SUM(add_fir[63:48]) );
  FIR_FILTER2_DW01_add_4 add_107 ( .A(fir_data[335:320]), .B(fir_data[191:176]), .SUM(add_fir[79:64]) );
  FIR_FILTER2_DW01_add_5 add_106 ( .A(fir_data[351:336]), .B(fir_data[175:160]), .SUM(add_fir[95:80]) );
  FIR_FILTER2_DW01_add_6 add_105 ( .A(fir_data[367:352]), .B(fir_data[159:144]), .SUM(add_fir[111:96]) );
  FIR_FILTER2_DW01_add_7 add_104 ( .A(fir_data[383:368]), .B(fir_data[143:128]), .SUM(add_fir[127:112]) );
  FIR_FILTER2_DW01_add_8 add_103 ( .A(fir_data[399:384]), .B(fir_data[127:112]), .SUM(add_fir[143:128]) );
  FIR_FILTER2_DW01_add_9 add_102 ( .A(fir_data[415:400]), .B(fir_data[111:96]), 
        .SUM(add_fir[159:144]) );
  FIR_FILTER2_DW01_add_10 add_101 ( .A(fir_data[431:416]), .B(fir_data[95:80]), 
        .SUM(add_fir[175:160]) );
  FIR_FILTER2_DW01_add_11 add_100 ( .A(fir_data[447:432]), .B(fir_data[79:64]), 
        .SUM(add_fir[191:176]) );
  FIR_FILTER2_DW01_add_12 add_99 ( .A(fir_data[463:448]), .B(fir_data[63:48]), 
        .SUM(add_fir[207:192]) );
  FIR_FILTER2_DW01_add_13 add_98 ( .A(fir_data[479:464]), .B(fir_data[47:32]), 
        .SUM(add_fir[223:208]) );
  FIR_FILTER2_DW01_add_14 add_97 ( .A(fir_data[495:480]), .B(fir_data[31:16]), 
        .SUM(add_fir[239:224]) );
  FIR_FILTER2_DW01_add_15 add_96 ( .A(fir_data[511:496]), .B(fir_data[15:0]), 
        .SUM(add_fir[255:240]) );
  FIR_FILTER2_DW01_add_30 add_172_12 ( .B(temp_mul_add_fir[31:0]), .SUM({N439, 
        N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, 
        N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, 
        N414, N413, N412, N411, N410, N409, N408}), .A_31_(
        temp_mul_add_fir[63]), .A_30_(temp_mul_add_fir[62]), .A_29_(
        temp_mul_add_fir[61]), .A_28_(temp_mul_add_fir[60]), .A_27_(
        temp_mul_add_fir[59]), .A_26_(temp_mul_add_fir[58]), .A_25_(
        temp_mul_add_fir[57]), .A_24_(temp_mul_add_fir[56]), .A_23_(
        temp_mul_add_fir[55]), .A_22_(temp_mul_add_fir[54]), .A_21_(
        temp_mul_add_fir[53]), .A_20_(temp_mul_add_fir[52]), .A_19_(
        temp_mul_add_fir[51]), .A_18_(temp_mul_add_fir[50]), .A_17_(
        temp_mul_add_fir[49]), .A_16_(temp_mul_add_fir[48]), .A_15_(
        temp_mul_add_fir[47]), .A_14_(temp_mul_add_fir[46]), .A_13_(
        temp_mul_add_fir[45]), .A_12_(temp_mul_add_fir[44]), .A_11_(
        temp_mul_add_fir[43]), .A_10_(temp_mul_add_fir[42]), .A_9_(
        temp_mul_add_fir[41]), .A_8_(temp_mul_add_fir[40]), .A_7_(
        temp_mul_add_fir[39]), .A_6_(temp_mul_add_fir[38]), .A_5_(
        temp_mul_add_fir[37]), .A_4_(temp_mul_add_fir[36]), .A_3_(
        temp_mul_add_fir[35]), .A_2_(temp_mul_add_fir[34]), .A_1_(
        temp_mul_add_fir[33]) );
  FIR_FILTER2_DW01_add_29 add_172_11 ( .A_31_(temp_mul_add_fir[127]), .A_30_(
        temp_mul_add_fir[126]), .A_29_(temp_mul_add_fir[125]), .A_28_(
        temp_mul_add_fir[124]), .A_27_(temp_mul_add_fir[123]), .A_26_(
        temp_mul_add_fir[122]), .A_25_(temp_mul_add_fir[121]), .A_24_(
        temp_mul_add_fir[120]), .A_23_(temp_mul_add_fir[119]), .A_22_(
        temp_mul_add_fir[118]), .A_21_(temp_mul_add_fir[117]), .A_20_(
        temp_mul_add_fir[116]), .A_19_(temp_mul_add_fir[115]), .A_18_(
        temp_mul_add_fir[114]), .A_17_(temp_mul_add_fir[113]), .A_16_(
        temp_mul_add_fir[112]), .A_15_(temp_mul_add_fir[111]), .A_14_(
        temp_mul_add_fir[110]), .A_13_(temp_mul_add_fir[109]), .A_12_(
        temp_mul_add_fir[108]), .A_11_(temp_mul_add_fir[107]), .A_10_(
        temp_mul_add_fir[106]), .A_9_(temp_mul_add_fir[105]), .A_8_(
        temp_mul_add_fir[104]), .A_7_(temp_mul_add_fir[103]), .A_6_(
        temp_mul_add_fir[102]), .A_5_(temp_mul_add_fir[101]), .A_4_(
        temp_mul_add_fir[100]), .A_3_(temp_mul_add_fir[99]), .A_2_(
        temp_mul_add_fir[98]), .A_1_(temp_mul_add_fir[97]), .B_31_(
        temp_mul_add_fir[95]), .B_30_(temp_mul_add_fir[94]), .B_29_(
        temp_mul_add_fir[93]), .B_28_(temp_mul_add_fir[92]), .B_27_(
        temp_mul_add_fir[91]), .B_26_(temp_mul_add_fir[90]), .B_25_(
        temp_mul_add_fir[89]), .B_24_(temp_mul_add_fir[88]), .B_23_(
        temp_mul_add_fir[87]), .B_22_(temp_mul_add_fir[86]), .B_21_(
        temp_mul_add_fir[85]), .B_20_(temp_mul_add_fir[84]), .B_19_(
        temp_mul_add_fir[83]), .B_18_(temp_mul_add_fir[82]), .B_17_(
        temp_mul_add_fir[81]), .B_16_(temp_mul_add_fir[80]), .B_15_(
        temp_mul_add_fir[79]), .B_14_(temp_mul_add_fir[78]), .B_13_(
        temp_mul_add_fir[77]), .B_12_(temp_mul_add_fir[76]), .B_11_(
        temp_mul_add_fir[75]), .B_10_(temp_mul_add_fir[74]), .B_9_(
        temp_mul_add_fir[73]), .B_8_(temp_mul_add_fir[72]), .B_7_(
        temp_mul_add_fir[71]), .B_6_(temp_mul_add_fir[70]), .B_5_(
        temp_mul_add_fir[69]), .B_4_(temp_mul_add_fir[68]), .B_3_(
        temp_mul_add_fir[67]), .B_2_(temp_mul_add_fir[66]), .SUM_31_(N407), 
        .SUM_30_(N406), .SUM_29_(N405), .SUM_28_(N404), .SUM_27_(N403), 
        .SUM_26_(N402), .SUM_25_(N401), .SUM_24_(N400), .SUM_23_(N399), 
        .SUM_22_(N398), .SUM_21_(N397), .SUM_20_(N396), .SUM_19_(N395), 
        .SUM_18_(N394), .SUM_17_(N393), .SUM_16_(N392), .SUM_15_(N391), 
        .SUM_14_(N390), .SUM_13_(N389), .SUM_12_(N388), .SUM_11_(N387), 
        .SUM_10_(N386), .SUM_9_(N385), .SUM_8_(N384), .SUM_7_(N383), .SUM_6_(
        N382), .SUM_5_(N381), .SUM_4_(N380), .SUM_3_(N379), .SUM_2_(N378), 
        .SUM_1_(N377) );
  FIR_FILTER2_DW01_add_28 add_172_9 ( .A_31_(temp_mul_add_fir[191]), .A_30_(
        temp_mul_add_fir[190]), .A_29_(temp_mul_add_fir[189]), .A_28_(
        temp_mul_add_fir[188]), .A_27_(temp_mul_add_fir[187]), .A_26_(
        temp_mul_add_fir[186]), .A_25_(temp_mul_add_fir[185]), .A_24_(
        temp_mul_add_fir[184]), .A_23_(temp_mul_add_fir[183]), .A_22_(
        temp_mul_add_fir[182]), .A_21_(temp_mul_add_fir[181]), .A_20_(
        temp_mul_add_fir[180]), .A_19_(temp_mul_add_fir[179]), .A_18_(
        temp_mul_add_fir[178]), .A_17_(temp_mul_add_fir[177]), .A_16_(
        temp_mul_add_fir[176]), .A_15_(temp_mul_add_fir[175]), .A_14_(
        temp_mul_add_fir[174]), .A_13_(temp_mul_add_fir[173]), .A_12_(
        temp_mul_add_fir[172]), .A_11_(temp_mul_add_fir[171]), .A_10_(
        temp_mul_add_fir[170]), .A_9_(temp_mul_add_fir[169]), .A_8_(
        temp_mul_add_fir[168]), .A_7_(temp_mul_add_fir[167]), .A_6_(
        temp_mul_add_fir[166]), .A_5_(temp_mul_add_fir[165]), .A_4_(
        temp_mul_add_fir[164]), .A_3_(temp_mul_add_fir[163]), .A_2_(
        temp_mul_add_fir[162]), .A_1_(temp_mul_add_fir[161]), .B_31_(
        temp_mul_add_fir[159]), .B_30_(temp_mul_add_fir[158]), .B_29_(
        temp_mul_add_fir[157]), .B_28_(temp_mul_add_fir[156]), .B_27_(
        temp_mul_add_fir[155]), .B_26_(temp_mul_add_fir[154]), .B_25_(
        temp_mul_add_fir[153]), .B_24_(temp_mul_add_fir[152]), .B_23_(
        temp_mul_add_fir[151]), .B_22_(temp_mul_add_fir[150]), .B_21_(
        temp_mul_add_fir[149]), .B_20_(temp_mul_add_fir[148]), .B_19_(
        temp_mul_add_fir[147]), .B_18_(temp_mul_add_fir[146]), .B_17_(
        temp_mul_add_fir[145]), .B_16_(temp_mul_add_fir[144]), .B_15_(
        temp_mul_add_fir[143]), .B_14_(temp_mul_add_fir[142]), .B_13_(
        temp_mul_add_fir[141]), .B_12_(temp_mul_add_fir[140]), .B_11_(
        temp_mul_add_fir[139]), .B_10_(temp_mul_add_fir[138]), .B_9_(
        temp_mul_add_fir[137]), .B_8_(temp_mul_add_fir[136]), .B_7_(
        temp_mul_add_fir[135]), .B_6_(temp_mul_add_fir[134]), .B_5_(
        temp_mul_add_fir[133]), .B_4_(temp_mul_add_fir[132]), .B_3_(
        temp_mul_add_fir[131]), .B_2_(temp_mul_add_fir[130]), .SUM_31_(N343), 
        .SUM_30_(N342), .SUM_29_(N341), .SUM_28_(N340), .SUM_27_(N339), 
        .SUM_26_(N338), .SUM_25_(N337), .SUM_24_(N336), .SUM_23_(N335), 
        .SUM_22_(N334), .SUM_21_(N333), .SUM_20_(N332), .SUM_19_(N331), 
        .SUM_18_(N330), .SUM_17_(N329), .SUM_16_(N328), .SUM_15_(N327), 
        .SUM_14_(N326), .SUM_13_(N325), .SUM_12_(N324), .SUM_11_(N323), 
        .SUM_10_(N322), .SUM_9_(N321), .SUM_8_(N320), .SUM_7_(N319), .SUM_6_(
        N318), .SUM_5_(N317), .SUM_4_(N316), .SUM_3_(N315), .SUM_2_(N314), 
        .SUM_1_(N313) );
  FIR_FILTER2_DW01_add_27 add_172_8 ( .A(temp_mul_add_fir[255:224]), .SUM({
        N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, 
        N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, 
        N287, N286, N285, N284, N283, N282, N281, N280}), .B_31_(
        temp_mul_add_fir[223]), .B_30_(temp_mul_add_fir[222]), .B_29_(
        temp_mul_add_fir[221]), .B_28_(temp_mul_add_fir[220]), .B_27_(
        temp_mul_add_fir[219]), .B_26_(temp_mul_add_fir[218]), .B_25_(
        temp_mul_add_fir[217]), .B_24_(temp_mul_add_fir[216]), .B_23_(
        temp_mul_add_fir[215]), .B_22_(temp_mul_add_fir[214]), .B_21_(
        temp_mul_add_fir[213]), .B_20_(temp_mul_add_fir[212]), .B_19_(
        temp_mul_add_fir[211]), .B_18_(temp_mul_add_fir[210]), .B_17_(
        temp_mul_add_fir[209]), .B_16_(temp_mul_add_fir[208]), .B_15_(
        temp_mul_add_fir[207]), .B_14_(temp_mul_add_fir[206]), .B_13_(
        temp_mul_add_fir[205]), .B_12_(temp_mul_add_fir[204]), .B_11_(
        temp_mul_add_fir[203]), .B_10_(temp_mul_add_fir[202]), .B_9_(
        temp_mul_add_fir[201]), .B_8_(temp_mul_add_fir[200]), .B_7_(
        temp_mul_add_fir[199]), .B_6_(temp_mul_add_fir[198]), .B_5_(
        temp_mul_add_fir[197]), .B_4_(temp_mul_add_fir[196]), .B_3_(
        temp_mul_add_fir[195]), .B_2_(temp_mul_add_fir[194]), .B_1_(
        temp_mul_add_fir[193]) );
  FIR_FILTER2_DW01_add_26 add_172_5 ( .A_31_(temp_mul_add_fir[319]), .A_30_(
        temp_mul_add_fir[318]), .A_29_(temp_mul_add_fir[317]), .A_28_(
        temp_mul_add_fir[316]), .A_27_(temp_mul_add_fir[315]), .A_26_(
        temp_mul_add_fir[314]), .A_25_(temp_mul_add_fir[313]), .A_24_(
        temp_mul_add_fir[312]), .A_23_(temp_mul_add_fir[311]), .A_22_(
        temp_mul_add_fir[310]), .A_21_(temp_mul_add_fir[309]), .A_20_(
        temp_mul_add_fir[308]), .A_19_(temp_mul_add_fir[307]), .A_18_(
        temp_mul_add_fir[306]), .A_17_(temp_mul_add_fir[305]), .A_16_(
        temp_mul_add_fir[304]), .A_15_(temp_mul_add_fir[303]), .A_14_(
        temp_mul_add_fir[302]), .A_13_(temp_mul_add_fir[301]), .A_12_(
        temp_mul_add_fir[300]), .A_11_(temp_mul_add_fir[299]), .A_10_(
        temp_mul_add_fir[298]), .A_9_(temp_mul_add_fir[297]), .A_8_(
        temp_mul_add_fir[296]), .A_7_(temp_mul_add_fir[295]), .A_6_(
        temp_mul_add_fir[294]), .A_5_(temp_mul_add_fir[293]), .A_4_(
        temp_mul_add_fir[292]), .A_3_(temp_mul_add_fir[291]), .A_2_(
        temp_mul_add_fir[290]), .A_1_(temp_mul_add_fir[289]), .B_31_(
        temp_mul_add_fir[287]), .B_30_(temp_mul_add_fir[286]), .B_29_(
        temp_mul_add_fir[285]), .B_28_(temp_mul_add_fir[284]), .B_27_(
        temp_mul_add_fir[283]), .B_26_(temp_mul_add_fir[282]), .B_25_(
        temp_mul_add_fir[281]), .B_24_(temp_mul_add_fir[280]), .B_23_(
        temp_mul_add_fir[279]), .B_22_(temp_mul_add_fir[278]), .B_21_(
        temp_mul_add_fir[277]), .B_20_(temp_mul_add_fir[276]), .B_19_(
        temp_mul_add_fir[275]), .B_18_(temp_mul_add_fir[274]), .B_17_(
        temp_mul_add_fir[273]), .B_16_(temp_mul_add_fir[272]), .B_15_(
        temp_mul_add_fir[271]), .B_14_(temp_mul_add_fir[270]), .B_13_(
        temp_mul_add_fir[269]), .B_12_(temp_mul_add_fir[268]), .B_11_(
        temp_mul_add_fir[267]), .B_10_(temp_mul_add_fir[266]), .B_9_(
        temp_mul_add_fir[265]), .B_8_(temp_mul_add_fir[264]), .B_7_(
        temp_mul_add_fir[263]), .B_6_(temp_mul_add_fir[262]), .B_5_(
        temp_mul_add_fir[261]), .B_4_(temp_mul_add_fir[260]), .B_3_(
        temp_mul_add_fir[259]), .B_2_(temp_mul_add_fir[258]), .SUM_31_(N215), 
        .SUM_30_(N214), .SUM_29_(N213), .SUM_28_(N212), .SUM_27_(N211), 
        .SUM_26_(N210), .SUM_25_(N209), .SUM_24_(N208), .SUM_23_(N207), 
        .SUM_22_(N206), .SUM_21_(N205), .SUM_20_(N204), .SUM_19_(N203), 
        .SUM_18_(N202), .SUM_17_(N201), .SUM_16_(N200), .SUM_15_(N199), 
        .SUM_14_(N198), .SUM_13_(N197), .SUM_12_(N196), .SUM_11_(N195), 
        .SUM_10_(N194), .SUM_9_(N193), .SUM_8_(N192), .SUM_7_(N191), .SUM_6_(
        N190), .SUM_5_(N189), .SUM_4_(N188), .SUM_3_(N187), .SUM_2_(N186), 
        .SUM_1_(N185) );
  FIR_FILTER2_DW01_add_25 add_172_4 ( .A(temp_mul_add_fir[383:352]), .SUM({
        N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, 
        N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, 
        N1600, N159, N158, N157, N156, N155, N154, N153, N152}), .B_31_(
        temp_mul_add_fir[351]), .B_30_(temp_mul_add_fir[350]), .B_29_(
        temp_mul_add_fir[349]), .B_28_(temp_mul_add_fir[348]), .B_27_(
        temp_mul_add_fir[347]), .B_26_(temp_mul_add_fir[346]), .B_25_(
        temp_mul_add_fir[345]), .B_24_(temp_mul_add_fir[344]), .B_23_(
        temp_mul_add_fir[343]), .B_22_(temp_mul_add_fir[342]), .B_21_(
        temp_mul_add_fir[341]), .B_20_(temp_mul_add_fir[340]), .B_19_(
        temp_mul_add_fir[339]), .B_18_(temp_mul_add_fir[338]), .B_17_(
        temp_mul_add_fir[337]), .B_16_(temp_mul_add_fir[336]), .B_15_(
        temp_mul_add_fir[335]), .B_14_(temp_mul_add_fir[334]), .B_13_(
        temp_mul_add_fir[333]), .B_12_(temp_mul_add_fir[332]), .B_11_(
        temp_mul_add_fir[331]), .B_10_(temp_mul_add_fir[330]), .B_9_(
        temp_mul_add_fir[329]), .B_8_(temp_mul_add_fir[328]), .B_7_(
        temp_mul_add_fir[327]), .B_6_(temp_mul_add_fir[326]), .B_5_(
        temp_mul_add_fir[325]), .B_4_(temp_mul_add_fir[324]), .B_3_(
        temp_mul_add_fir[323]), .B_2_(temp_mul_add_fir[322]), .B_1_(
        temp_mul_add_fir[321]) );
  FIR_FILTER2_DW01_add_24 add_172_2 ( .A(temp_mul_add_fir[447:416]), .B(
        temp_mul_add_fir[415:384]), .SUM({N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88}) );
  FIR_FILTER2_DW01_add_23 add_172 ( .A_31_(temp_mul_add_fir[511]), .A_30_(
        temp_mul_add_fir[510]), .A_29_(temp_mul_add_fir[509]), .A_28_(
        temp_mul_add_fir[508]), .A_27_(temp_mul_add_fir[507]), .A_26_(
        temp_mul_add_fir[506]), .A_25_(temp_mul_add_fir[505]), .A_24_(
        temp_mul_add_fir[504]), .A_23_(temp_mul_add_fir[503]), .A_22_(
        temp_mul_add_fir[502]), .A_21_(temp_mul_add_fir[501]), .A_20_(
        temp_mul_add_fir[500]), .A_19_(temp_mul_add_fir[499]), .A_18_(
        temp_mul_add_fir[498]), .A_17_(temp_mul_add_fir[497]), .A_16_(
        temp_mul_add_fir[496]), .A_15_(temp_mul_add_fir[495]), .A_14_(
        temp_mul_add_fir[494]), .A_13_(temp_mul_add_fir[493]), .A_12_(
        temp_mul_add_fir[492]), .A_11_(temp_mul_add_fir[491]), .A_10_(
        temp_mul_add_fir[490]), .A_9_(temp_mul_add_fir[489]), .A_8_(
        temp_mul_add_fir[488]), .A_7_(temp_mul_add_fir[487]), .A_6_(
        temp_mul_add_fir[486]), .A_5_(temp_mul_add_fir[485]), .A_4_(
        temp_mul_add_fir[484]), .A_3_(temp_mul_add_fir[483]), .A_2_(
        temp_mul_add_fir[482]), .A_1_(temp_mul_add_fir[481]), .B_31_(
        temp_mul_add_fir[479]), .B_30_(temp_mul_add_fir[478]), .B_29_(
        temp_mul_add_fir[477]), .B_28_(temp_mul_add_fir[476]), .B_27_(
        temp_mul_add_fir[475]), .B_26_(temp_mul_add_fir[474]), .B_25_(
        temp_mul_add_fir[473]), .B_24_(temp_mul_add_fir[472]), .B_23_(
        temp_mul_add_fir[471]), .B_22_(temp_mul_add_fir[470]), .B_21_(
        temp_mul_add_fir[469]), .B_20_(temp_mul_add_fir[468]), .B_19_(
        temp_mul_add_fir[467]), .B_18_(temp_mul_add_fir[466]), .B_17_(
        temp_mul_add_fir[465]), .B_16_(temp_mul_add_fir[464]), .B_15_(
        temp_mul_add_fir[463]), .B_14_(temp_mul_add_fir[462]), .B_13_(
        temp_mul_add_fir[461]), .B_12_(temp_mul_add_fir[460]), .B_11_(
        temp_mul_add_fir[459]), .B_10_(temp_mul_add_fir[458]), .B_9_(
        temp_mul_add_fir[457]), .B_8_(temp_mul_add_fir[456]), .B_7_(
        temp_mul_add_fir[455]), .B_6_(temp_mul_add_fir[454]), .B_5_(
        temp_mul_add_fir[453]), .B_4_(temp_mul_add_fir[452]), .B_3_(
        temp_mul_add_fir[451]), .B_2_(temp_mul_add_fir[450]), .B_1_(
        temp_mul_add_fir[449]), .SUM_31_(N87), .SUM_30_(N86), .SUM_29_(N85), 
        .SUM_28_(N84), .SUM_27_(N83), .SUM_26_(N82), .SUM_25_(N81), .SUM_24_(
        N80), .SUM_23_(N79), .SUM_22_(N78), .SUM_21_(N77), .SUM_20_(N76), 
        .SUM_19_(N75), .SUM_18_(N74), .SUM_17_(N73), .SUM_16_(N720), .SUM_15_(
        N710), .SUM_14_(N702), .SUM_13_(N690), .SUM_12_(N680), .SUM_11_(N670), 
        .SUM_10_(N660), .SUM_9_(N650), .SUM_8_(N640), .SUM_7_(N630), .SUM_6_(
        N620), .SUM_5_(N610), .SUM_4_(N600), .SUM_3_(N590), .SUM_2_(N580), 
        .SUM_1_(N57) );
  FIR_FILTER2_DW01_add_22 add_172_13 ( .B({N439, N438, N437, N436, N435, N434, 
        N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, 
        N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, 
        N409, N408}), .SUM({N471, N470, N469, N468, N467, N466, N465, N464, 
        N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, 
        N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440}), .A_31_(N407), .A_30_(N406), .A_29_(N405), .A_28_(N404), .A_27_(N403), 
        .A_26_(N402), .A_25_(N401), .A_24_(N400), .A_23_(N399), .A_22_(N398), 
        .A_21_(N397), .A_20_(N396), .A_19_(N395), .A_18_(N394), .A_17_(N393), 
        .A_16_(N392), .A_15_(N391), .A_14_(N390), .A_13_(N389), .A_12_(N388), 
        .A_11_(N387), .A_10_(N386), .A_9_(N385), .A_8_(N384), .A_7_(N383), 
        .A_6_(N382), .A_5_(N381), .A_4_(N380), .A_3_(N379), .A_2_(N378), 
        .A_1_(N377) );
  FIR_FILTER2_DW01_add_21 add_172_10 ( .A({N311, N310, N309, N308, N307, N306, 
        N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, 
        N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280}), .SUM({N375, N374, N373, N372, N371, N370, N369, N368, 
        N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, 
        N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344}), .B_31_(N343), .B_30_(N342), .B_29_(N341), .B_28_(N340), .B_27_(N339), 
        .B_26_(N338), .B_25_(N337), .B_24_(N336), .B_23_(N335), .B_22_(N334), 
        .B_21_(N333), .B_20_(N332), .B_19_(N331), .B_18_(N330), .B_17_(N329), 
        .B_16_(N328), .B_15_(N327), .B_14_(N326), .B_13_(N325), .B_12_(N324), 
        .B_11_(N323), .B_10_(N322), .B_9_(N321), .B_8_(N320), .B_7_(N319), 
        .B_6_(N318), .B_5_(N317), .B_4_(N316), .B_3_(N315), .B_2_(N314), 
        .B_1_(N313) );
  FIR_FILTER2_DW01_add_20 add_172_6 ( .A({N183, N182, N181, N180, N179, N178, 
        N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, 
        N165, N164, N163, N162, N161, N1600, N159, N158, N157, N156, N155, 
        N154, N153, N152}), .SUM({N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216}), .B_31_(N215), .B_30_(N214), .B_29_(N213), .B_28_(N212), 
        .B_27_(N211), .B_26_(N210), .B_25_(N209), .B_24_(N208), .B_23_(N207), 
        .B_22_(N206), .B_21_(N205), .B_20_(N204), .B_19_(N203), .B_18_(N202), 
        .B_17_(N201), .B_16_(N200), .B_15_(N199), .B_14_(N198), .B_13_(N197), 
        .B_12_(N196), .B_11_(N195), .B_10_(N194), .B_9_(N193), .B_8_(N192), 
        .B_7_(N191), .B_6_(N190), .B_5_(N189), .B_4_(N188), .B_3_(N187), 
        .B_2_(N186), .B_1_(N185) );
  FIR_FILTER2_DW01_add_19 add_172_3 ( .B({N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88}), .SUM({N151, N1500, N1490, N148, N147, N146, N145, N144, N143, N142, N141, 
        N1401, N139, N138, N137, N136, N135, N134, N133, N132, N131, N1301, 
        N129, N128, N127, N126, N125, N124, N123, N122, N121, N1201}), .A_31_(
        N87), .A_30_(N86), .A_29_(N85), .A_28_(N84), .A_27_(N83), .A_26_(N82), 
        .A_25_(N81), .A_24_(N80), .A_23_(N79), .A_22_(N78), .A_21_(N77), 
        .A_20_(N76), .A_19_(N75), .A_18_(N74), .A_17_(N73), .A_16_(N720), 
        .A_15_(N710), .A_14_(N702), .A_13_(N690), .A_12_(N680), .A_11_(N670), 
        .A_10_(N660), .A_9_(N650), .A_8_(N640), .A_7_(N630), .A_6_(N620), 
        .A_5_(N610), .A_4_(N600), .A_3_(N590), .A_2_(N580), .A_1_(N57) );
  FIR_FILTER2_DW01_add_18 add_172_14 ( .A({N375, N374, N373, N372, N371, N370, 
        N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, 
        N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, 
        N345, N344}), .B({N471, N470, N469, N468, N467, N466, N465, N464, N463, 
        N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, 
        N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440}), 
        .SUM({N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, 
        N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, 
        N480, N479, N478, N477, N476, N475, N474, N473, N472}) );
  FIR_FILTER2_DW01_add_17 add_172_7 ( .A({N151, N1500, N1490, N148, N147, N146, 
        N145, N144, N143, N142, N141, N1401, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N1301, N129, N128, N127, N126, N125, N124, 
        N123, N122, N121, N1201}), .B({N247, N246, N245, N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, 
        N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, 
        N217, N216}), .SUM({N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248}) );
  FIR_FILTER2_DW01_add_16 add_172_15 ( .A({N279, N278, N277, N276, N275, N274, 
        N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, 
        N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, 
        N249, N248}), .B({N503, N502, N501, N500, N499, N498, N497, N496, N495, 
        N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, 
        N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472}), 
        .SUM_31_(comb_fir_o[31]), .SUM_30_(comb_fir_o[30]), .SUM_29_(
        comb_fir_o[29]), .SUM_28_(comb_fir_o[28]), .SUM_27_(comb_fir_o[27]), 
        .SUM_26_(comb_fir_o[26]), .SUM_25_(comb_fir_o[25]), .SUM_24_(
        comb_fir_o[24]), .SUM_23_(comb_fir_o[23]), .SUM_22_(comb_fir_o[22]), 
        .SUM_21_(comb_fir_o[21]), .SUM_20_(comb_fir_o[20]), .SUM_19_(
        comb_fir_o[19]), .SUM_18_(comb_fir_o[18]), .SUM_17_(comb_fir_o[17]), 
        .SUM_16_(comb_fir_o[16]) );
  FIR_FILTER2_DW01_inc_1 add_177 ( .A({n540, comb_fir_o[30:16]}), .SUM({N520, 
        N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, 
        N507, N506, N505}) );
  FIR_FILTER2_DW_mult_uns_15 mult_113 ( .a_15_(temp_add_fir[252]), .a_14_(
        temp_add_fir[251]), .a_13_(temp_add_fir[250]), .a_12_(
        temp_add_fir[249]), .a_11_(temp_add_fir[248]), .a_10_(
        temp_add_fir[247]), .a_9_(temp_add_fir[246]), .a_8_(temp_add_fir[245]), 
        .a_7_(temp_add_fir[244]), .a_6_(temp_add_fir[243]), .a_5_(
        temp_add_fir[242]), .a_4_(temp_add_fir[241]), .a_3_(temp_add_fir[240]), 
        .a_2_(temp_add_fir[239]), .a_1_(temp_add_fir[238]), .a_0_(
        temp_add_fir[237]), .product_31_(mul_add_fir[487]), .product_30_(
        mul_add_fir[486]), .product_29_(mul_add_fir[485]), .product_28_(
        mul_add_fir[484]), .product_27_(mul_add_fir[483]), .product_26_(
        mul_add_fir[482]), .product_25_(mul_add_fir[481]), .product_24_(
        mul_add_fir[480]), .product_23_(mul_add_fir[479]), .product_22_(
        mul_add_fir[478]), .product_21_(mul_add_fir[477]), .product_20_(
        mul_add_fir[476]), .product_19_(mul_add_fir[475]), .product_18_(
        mul_add_fir[474]), .product_17_(mul_add_fir[473]), .product_16_(
        mul_add_fir[472]), .product_15_(mul_add_fir[471]), .product_14_(
        mul_add_fir[470]), .product_13_(mul_add_fir[469]), .product_12_(
        mul_add_fir[468]), .product_11_(mul_add_fir[467]), .product_10_(
        mul_add_fir[466]), .product_9_(mul_add_fir[465]), .product_8_(
        mul_add_fir[464]), .product_7_(mul_add_fir[463]), .product_6_(
        mul_add_fir[462]), .product_5_(mul_add_fir[461]), .product_4_(
        mul_add_fir[460]), .product_3_(mul_add_fir[459]), .product_2_(
        mul_add_fir[458]), .product_1_(mul_add_fir[457]) );
  FIR_FILTER2_DW_mult_uns_14 mult_114 ( .a_15_(temp_add_fir[236]), .a_14_(
        temp_add_fir[235]), .a_13_(temp_add_fir[234]), .a_12_(
        temp_add_fir[233]), .a_11_(temp_add_fir[232]), .a_10_(
        temp_add_fir[231]), .a_9_(temp_add_fir[230]), .a_8_(temp_add_fir[229]), 
        .a_7_(temp_add_fir[228]), .a_6_(temp_add_fir[227]), .a_5_(
        temp_add_fir[226]), .a_4_(temp_add_fir[225]), .a_3_(temp_add_fir[224]), 
        .a_2_(temp_add_fir[223]), .a_1_(temp_add_fir[222]), .a_0_(
        temp_add_fir[221]), .product_31_(mul_add_fir[456]), .product_30_(
        mul_add_fir[455]), .product_29_(mul_add_fir[454]), .product_28_(
        mul_add_fir[453]), .product_27_(mul_add_fir[452]), .product_26_(
        mul_add_fir[451]), .product_25_(mul_add_fir[450]), .product_24_(
        mul_add_fir[449]), .product_23_(mul_add_fir[448]), .product_22_(
        mul_add_fir[447]), .product_21_(mul_add_fir[446]), .product_20_(
        mul_add_fir[445]), .product_19_(mul_add_fir[444]), .product_18_(
        mul_add_fir[443]), .product_17_(mul_add_fir[442]), .product_16_(
        mul_add_fir[441]), .product_15_(mul_add_fir[440]), .product_14_(
        mul_add_fir[439]), .product_13_(mul_add_fir[438]), .product_12_(
        mul_add_fir[437]), .product_11_(mul_add_fir[436]), .product_10_(
        mul_add_fir[435]), .product_9_(mul_add_fir[434]), .product_8_(
        mul_add_fir[433]), .product_7_(mul_add_fir[432]), .product_6_(
        mul_add_fir[431]), .product_5_(mul_add_fir[430]), .product_4_(
        mul_add_fir[429]), .product_3_(mul_add_fir[428]), .product_2_(
        mul_add_fir[427]), .product_1_(mul_add_fir[426]) );
  FIR_FILTER2_DW_mult_uns_13 mult_115 ( .a_15_(temp_add_fir[220]), .a_14_(
        temp_add_fir[219]), .a_13_(temp_add_fir[218]), .a_12_(
        temp_add_fir[217]), .a_11_(temp_add_fir[216]), .a_10_(
        temp_add_fir[215]), .a_9_(temp_add_fir[214]), .a_8_(temp_add_fir[213]), 
        .a_7_(temp_add_fir[212]), .a_6_(temp_add_fir[211]), .a_5_(
        temp_add_fir[210]), .a_4_(temp_add_fir[209]), .a_3_(temp_add_fir[208]), 
        .a_2_(temp_add_fir[207]), .a_1_(temp_add_fir[206]), .a_0_(
        temp_add_fir[205]), .product_31_(mul_add_fir[425]), .product_30_(
        mul_add_fir[424]), .product_29_(mul_add_fir[423]), .product_28_(
        mul_add_fir[422]), .product_27_(mul_add_fir[421]), .product_26_(
        mul_add_fir[420]), .product_25_(mul_add_fir[419]), .product_24_(
        mul_add_fir[418]), .product_23_(mul_add_fir[417]), .product_22_(
        mul_add_fir[416]), .product_21_(mul_add_fir[415]), .product_20_(
        mul_add_fir[414]), .product_19_(mul_add_fir[413]), .product_18_(
        mul_add_fir[412]), .product_17_(mul_add_fir[411]), .product_16_(
        mul_add_fir[410]), .product_15_(mul_add_fir[409]), .product_14_(
        mul_add_fir[408]), .product_13_(mul_add_fir[407]), .product_12_(
        mul_add_fir[406]), .product_11_(mul_add_fir[405]), .product_10_(
        mul_add_fir[404]), .product_9_(mul_add_fir[403]), .product_8_(
        mul_add_fir[402]), .product_7_(mul_add_fir[401]), .product_6_(
        mul_add_fir[400]), .product_5_(mul_add_fir[399]), .product_4_(
        mul_add_fir[398]), .product_3_(mul_add_fir[397]), .product_2_(
        mul_add_fir[396]), .product_1_(mul_add_fir[395]), .product_0_(
        mul_add_fir[394]) );
  FIR_FILTER2_DW_mult_uns_12 mult_116 ( .a_15_(temp_add_fir[204]), .a_14_(
        temp_add_fir[203]), .a_13_(temp_add_fir[202]), .a_12_(
        temp_add_fir[201]), .a_11_(temp_add_fir[200]), .a_10_(
        temp_add_fir[199]), .a_9_(temp_add_fir[198]), .a_8_(temp_add_fir[197]), 
        .a_7_(temp_add_fir[196]), .a_6_(temp_add_fir[195]), .a_5_(
        temp_add_fir[194]), .a_4_(temp_add_fir[193]), .a_3_(temp_add_fir[192]), 
        .a_2_(temp_add_fir[191]), .a_1_(temp_add_fir[190]), .a_0_(
        temp_add_fir[189]), .product_31_(mul_add_fir[393]), .product_30_(
        mul_add_fir[392]), .product_29_(mul_add_fir[391]), .product_28_(
        mul_add_fir[390]), .product_27_(mul_add_fir[389]), .product_26_(
        mul_add_fir[388]), .product_25_(mul_add_fir[387]), .product_24_(
        mul_add_fir[386]), .product_23_(mul_add_fir[385]), .product_22_(
        mul_add_fir[384]), .product_21_(mul_add_fir[383]), .product_20_(
        mul_add_fir[382]), .product_19_(mul_add_fir[381]), .product_18_(
        mul_add_fir[380]), .product_17_(mul_add_fir[379]), .product_16_(
        mul_add_fir[378]), .product_15_(mul_add_fir[377]), .product_14_(
        mul_add_fir[376]), .product_13_(mul_add_fir[375]), .product_12_(
        mul_add_fir[374]), .product_11_(mul_add_fir[373]), .product_10_(
        mul_add_fir[372]), .product_9_(mul_add_fir[371]), .product_8_(
        mul_add_fir[370]), .product_7_(mul_add_fir[369]), .product_6_(
        mul_add_fir[368]), .product_5_(mul_add_fir[367]), .product_4_(
        mul_add_fir[366]), .product_3_(mul_add_fir[365]), .product_2_(
        mul_add_fir[364]), .product_1_(mul_add_fir[363]), .product_0_(
        mul_add_fir[362]) );
  FIR_FILTER2_DW_mult_uns_11 mult_117 ( .a_16_(temp_add_fir[188]), .a_15_(
        temp_add_fir[188]), .a_14_(temp_add_fir[187]), .a_13_(
        temp_add_fir[186]), .a_12_(temp_add_fir[185]), .a_11_(
        temp_add_fir[184]), .a_10_(temp_add_fir[183]), .a_9_(temp_add_fir[182]), .a_8_(temp_add_fir[181]), .a_7_(temp_add_fir[180]), .a_6_(temp_add_fir[179]), 
        .a_5_(temp_add_fir[178]), .a_4_(temp_add_fir[177]), .a_3_(
        temp_add_fir[176]), .a_2_(temp_add_fir[175]), .a_1_(temp_add_fir[174]), 
        .a_0_(temp_add_fir[173]), .product_31_(mul_add_fir[361]), 
        .product_30_(mul_add_fir[360]), .product_29_(mul_add_fir[359]), 
        .product_28_(mul_add_fir[358]), .product_27_(mul_add_fir[357]), 
        .product_26_(mul_add_fir[356]), .product_25_(mul_add_fir[355]), 
        .product_24_(mul_add_fir[354]), .product_23_(mul_add_fir[353]), 
        .product_22_(mul_add_fir[352]), .product_21_(mul_add_fir[351]), 
        .product_20_(mul_add_fir[350]), .product_19_(mul_add_fir[349]), 
        .product_18_(mul_add_fir[348]), .product_17_(mul_add_fir[347]), 
        .product_16_(mul_add_fir[346]), .product_15_(mul_add_fir[345]), 
        .product_14_(mul_add_fir[344]), .product_13_(mul_add_fir[343]), 
        .product_12_(mul_add_fir[342]), .product_11_(mul_add_fir[341]), 
        .product_10_(mul_add_fir[340]), .product_9_(mul_add_fir[339]), 
        .product_8_(mul_add_fir[338]), .product_7_(mul_add_fir[337]), 
        .product_6_(mul_add_fir[336]), .product_5_(mul_add_fir[335]), 
        .product_4_(mul_add_fir[334]), .product_3_(mul_add_fir[333]), 
        .product_2_(mul_add_fir[332]), .product_1_(mul_add_fir[331]), 
        .product_0_(mul_add_fir[330]) );
  FIR_FILTER2_DW_mult_uns_10 mult_118 ( .a_16_(n740), .a_15_(n740), .a_14_(
        temp_add_fir[171]), .a_13_(temp_add_fir[170]), .a_12_(
        temp_add_fir[169]), .a_11_(temp_add_fir[168]), .a_10_(
        temp_add_fir[167]), .a_9_(temp_add_fir[166]), .a_8_(temp_add_fir[165]), 
        .a_7_(temp_add_fir[164]), .a_6_(temp_add_fir[163]), .a_5_(
        temp_add_fir[162]), .a_4_(temp_add_fir[161]), .a_3_(temp_add_fir[160]), 
        .a_2_(temp_add_fir[159]), .a_1_(temp_add_fir[158]), .a_0_(
        temp_add_fir[157]), .product_31_(mul_add_fir[329]), .product_30_(
        mul_add_fir[328]), .product_29_(mul_add_fir[327]), .product_28_(
        mul_add_fir[326]), .product_27_(mul_add_fir[325]), .product_26_(
        mul_add_fir[324]), .product_25_(mul_add_fir[323]), .product_24_(
        mul_add_fir[322]), .product_23_(mul_add_fir[321]), .product_22_(
        mul_add_fir[320]), .product_21_(mul_add_fir[319]), .product_20_(
        mul_add_fir[318]), .product_19_(mul_add_fir[317]), .product_18_(
        mul_add_fir[316]), .product_17_(mul_add_fir[315]), .product_16_(
        mul_add_fir[314]), .product_15_(mul_add_fir[313]), .product_14_(
        mul_add_fir[312]), .product_13_(mul_add_fir[311]), .product_12_(
        mul_add_fir[310]), .product_11_(mul_add_fir[309]), .product_10_(
        mul_add_fir[308]), .product_9_(mul_add_fir[307]), .product_8_(
        mul_add_fir[306]), .product_7_(mul_add_fir[305]), .product_6_(
        mul_add_fir[304]), .product_5_(mul_add_fir[303]), .product_4_(
        mul_add_fir[302]), .product_3_(mul_add_fir[301]), .product_2_(
        mul_add_fir[300]), .product_1_(mul_add_fir[299]) );
  FIR_FILTER2_DW_mult_uns_9 mult_119 ( .a_16_(n730), .a_15_(n730), .a_14_(
        temp_add_fir[155]), .a_13_(temp_add_fir[154]), .a_12_(
        temp_add_fir[153]), .a_11_(temp_add_fir[152]), .a_10_(
        temp_add_fir[151]), .a_9_(temp_add_fir[150]), .a_8_(temp_add_fir[149]), 
        .a_7_(temp_add_fir[148]), .a_6_(temp_add_fir[147]), .a_5_(
        temp_add_fir[146]), .a_4_(temp_add_fir[145]), .a_3_(temp_add_fir[144]), 
        .a_2_(temp_add_fir[143]), .a_1_(temp_add_fir[142]), .a_0_(
        temp_add_fir[141]), .product_31_(mul_add_fir[298]), .product_30_(
        mul_add_fir[297]), .product_29_(mul_add_fir[296]), .product_28_(
        mul_add_fir[295]), .product_27_(mul_add_fir[294]), .product_26_(
        mul_add_fir[293]), .product_25_(mul_add_fir[292]), .product_24_(
        mul_add_fir[291]), .product_23_(mul_add_fir[290]), .product_22_(
        mul_add_fir[289]), .product_21_(mul_add_fir[288]), .product_20_(
        mul_add_fir[287]), .product_19_(mul_add_fir[286]), .product_18_(
        mul_add_fir[285]), .product_17_(mul_add_fir[284]), .product_16_(
        mul_add_fir[283]), .product_15_(mul_add_fir[282]), .product_14_(
        mul_add_fir[281]), .product_13_(mul_add_fir[280]), .product_12_(
        mul_add_fir[279]), .product_11_(mul_add_fir[278]), .product_10_(
        mul_add_fir[277]), .product_9_(mul_add_fir[276]), .product_8_(
        mul_add_fir[275]), .product_7_(mul_add_fir[274]), .product_6_(
        mul_add_fir[273]), .product_5_(mul_add_fir[272]), .product_4_(
        mul_add_fir[271]), .product_3_(mul_add_fir[270]), .product_2_(
        mul_add_fir[269]), .product_1_(mul_add_fir[268]) );
  FIR_FILTER2_DW_mult_uns_7 mult_121 ( .a_15_(temp_add_fir[127]), .a_14_(
        temp_add_fir[126]), .a_13_(temp_add_fir[125]), .a_12_(
        temp_add_fir[124]), .a_11_(temp_add_fir[123]), .a_10_(
        temp_add_fir[122]), .a_9_(temp_add_fir[121]), .a_8_(temp_add_fir[120]), 
        .a_7_(temp_add_fir[119]), .a_6_(temp_add_fir[118]), .a_5_(
        temp_add_fir[117]), .a_4_(temp_add_fir[116]), .a_3_(temp_add_fir[115]), 
        .a_2_(temp_add_fir[114]), .a_1_(temp_add_fir[113]), .a_0_(
        temp_add_fir[112]), .product_31_(mul_add_fir[247]), .product_30_(
        mul_add_fir[246]), .product_29_(mul_add_fir[245]), .product_28_(
        mul_add_fir[244]), .product_27_(mul_add_fir[243]), .product_26_(
        mul_add_fir[242]), .product_25_(mul_add_fir[241]), .product_24_(
        mul_add_fir[240]), .product_23_(mul_add_fir[239]), .product_22_(
        mul_add_fir[238]), .product_21_(mul_add_fir[237]), .product_20_(
        mul_add_fir[236]), .product_19_(mul_add_fir[235]), .product_18_(
        mul_add_fir[234]), .product_17_(mul_add_fir[233]), .product_16_(
        mul_add_fir[232]), .product_15_(mul_add_fir[231]), .product_14_(
        mul_add_fir[230]), .product_13_(mul_add_fir[229]), .product_12_(
        mul_add_fir[228]), .product_11_(mul_add_fir[227]), .product_10_(
        mul_add_fir[226]), .product_9_(mul_add_fir[225]), .product_8_(
        mul_add_fir[224]), .product_7_(mul_add_fir[223]), .product_6_(
        mul_add_fir[222]), .product_5_(mul_add_fir[221]), .product_4_(
        mul_add_fir[220]), .product_3_(mul_add_fir[219]), .product_2_(
        mul_add_fir[218]), .product_1_(mul_add_fir[217]), .product_0_(
        mul_add_fir[216]) );
  FIR_FILTER2_DW_mult_uns_6 mult_122 ( .a_15_(temp_add_fir[111]), .a_14_(
        temp_add_fir[110]), .a_13_(temp_add_fir[109]), .a_12_(
        temp_add_fir[108]), .a_11_(temp_add_fir[107]), .a_10_(
        temp_add_fir[106]), .a_9_(temp_add_fir[105]), .a_8_(temp_add_fir[104]), 
        .a_7_(temp_add_fir[103]), .a_6_(temp_add_fir[102]), .a_5_(
        temp_add_fir[101]), .a_4_(temp_add_fir[100]), .a_3_(temp_add_fir[99]), 
        .a_2_(temp_add_fir[98]), .a_1_(temp_add_fir[97]), .a_0_(
        temp_add_fir[96]), .product_31_(mul_add_fir[215]), .product_30_(
        mul_add_fir[214]), .product_29_(mul_add_fir[213]), .product_28_(
        mul_add_fir[212]), .product_27_(mul_add_fir[211]), .product_26_(
        mul_add_fir[210]), .product_25_(mul_add_fir[209]), .product_24_(
        mul_add_fir[208]), .product_23_(mul_add_fir[207]), .product_22_(
        mul_add_fir[206]), .product_21_(mul_add_fir[205]), .product_20_(
        mul_add_fir[204]), .product_19_(mul_add_fir[203]), .product_18_(
        mul_add_fir[202]), .product_17_(mul_add_fir[201]), .product_16_(
        mul_add_fir[200]), .product_15_(mul_add_fir[199]), .product_14_(
        mul_add_fir[198]), .product_13_(mul_add_fir[197]), .product_12_(
        mul_add_fir[196]), .product_11_(mul_add_fir[195]), .product_10_(
        mul_add_fir[194]), .product_9_(mul_add_fir[193]), .product_8_(
        mul_add_fir[192]), .product_7_(mul_add_fir[191]), .product_6_(
        mul_add_fir[190]), .product_5_(mul_add_fir[189]), .product_4_(
        mul_add_fir[188]), .product_3_(mul_add_fir[187]), .product_2_(
        mul_add_fir[186]), .product_1_(mul_add_fir[185]) );
  FIR_FILTER2_DW_mult_uns_5 mult_123 ( .a_15_(temp_add_fir[95]), .a_14_(
        temp_add_fir[94]), .a_13_(temp_add_fir[93]), .a_12_(temp_add_fir[92]), 
        .a_11_(temp_add_fir[91]), .a_10_(temp_add_fir[90]), .a_9_(
        temp_add_fir[89]), .a_8_(temp_add_fir[88]), .a_7_(temp_add_fir[87]), 
        .a_6_(temp_add_fir[86]), .a_5_(temp_add_fir[85]), .a_4_(
        temp_add_fir[84]), .a_3_(temp_add_fir[83]), .a_2_(temp_add_fir[82]), 
        .a_1_(temp_add_fir[81]), .a_0_(temp_add_fir[80]), .product_31_(
        mul_add_fir[184]), .product_30_(mul_add_fir[183]), .product_29_(
        mul_add_fir[182]), .product_28_(mul_add_fir[181]), .product_27_(
        mul_add_fir[180]), .product_26_(mul_add_fir[179]), .product_25_(
        mul_add_fir[178]), .product_24_(mul_add_fir[177]), .product_23_(
        mul_add_fir[176]), .product_22_(mul_add_fir[175]), .product_21_(
        mul_add_fir[174]), .product_20_(mul_add_fir[173]), .product_19_(
        mul_add_fir[172]), .product_18_(mul_add_fir[171]), .product_17_(
        mul_add_fir[170]), .product_16_(mul_add_fir[169]), .product_15_(
        mul_add_fir[168]), .product_14_(mul_add_fir[167]), .product_13_(
        mul_add_fir[166]), .product_12_(mul_add_fir[165]), .product_11_(
        mul_add_fir[164]), .product_10_(mul_add_fir[163]), .product_9_(
        mul_add_fir[162]), .product_8_(mul_add_fir[161]), .product_7_(
        mul_add_fir[160]), .product_6_(mul_add_fir[159]), .product_5_(
        mul_add_fir[158]), .product_4_(mul_add_fir[157]), .product_3_(
        mul_add_fir[156]), .product_2_(mul_add_fir[155]), .product_1_(
        mul_add_fir[154]) );
  FIR_FILTER2_DW_mult_uns_4 mult_124 ( .a_16_(temp_add_fir[79]), .a_15_(
        temp_add_fir[79]), .a_14_(temp_add_fir[78]), .a_13_(temp_add_fir[77]), 
        .a_12_(temp_add_fir[76]), .a_11_(temp_add_fir[75]), .a_10_(
        temp_add_fir[74]), .a_9_(temp_add_fir[73]), .a_8_(temp_add_fir[72]), 
        .a_7_(temp_add_fir[71]), .a_6_(temp_add_fir[70]), .a_5_(
        temp_add_fir[69]), .a_4_(temp_add_fir[68]), .a_3_(temp_add_fir[67]), 
        .a_2_(temp_add_fir[66]), .a_1_(temp_add_fir[65]), .a_0_(
        temp_add_fir[64]), .product_31_(mul_add_fir[153]), .product_30_(
        mul_add_fir[152]), .product_29_(mul_add_fir[151]), .product_28_(
        mul_add_fir[150]), .product_27_(mul_add_fir[149]), .product_26_(
        mul_add_fir[148]), .product_25_(mul_add_fir[147]), .product_24_(
        mul_add_fir[146]), .product_23_(mul_add_fir[145]), .product_22_(
        mul_add_fir[144]), .product_21_(mul_add_fir[143]), .product_20_(
        mul_add_fir[142]), .product_19_(mul_add_fir[141]), .product_18_(
        mul_add_fir[140]), .product_17_(mul_add_fir[139]), .product_16_(
        mul_add_fir[138]), .product_15_(mul_add_fir[137]), .product_14_(
        mul_add_fir[136]), .product_13_(mul_add_fir[135]), .product_12_(
        mul_add_fir[134]), .product_11_(mul_add_fir[133]), .product_10_(
        mul_add_fir[132]), .product_9_(mul_add_fir[131]), .product_8_(
        mul_add_fir[130]), .product_7_(mul_add_fir[129]), .product_6_(
        mul_add_fir[128]), .product_5_(mul_add_fir[127]), .product_4_(
        mul_add_fir[126]), .product_3_(mul_add_fir[125]), .product_2_(
        mul_add_fir[124]) );
  FIR_FILTER2_DW_mult_uns_3 mult_125 ( .a_16_(n570), .a_15_(n570), .a_14_(
        temp_add_fir[62]), .a_13_(temp_add_fir[61]), .a_12_(temp_add_fir[60]), 
        .a_11_(temp_add_fir[59]), .a_10_(temp_add_fir[58]), .a_9_(
        temp_add_fir[57]), .a_8_(temp_add_fir[56]), .a_7_(temp_add_fir[55]), 
        .a_6_(temp_add_fir[54]), .a_5_(temp_add_fir[53]), .a_4_(
        temp_add_fir[52]), .a_3_(temp_add_fir[51]), .a_2_(temp_add_fir[50]), 
        .a_1_(temp_add_fir[49]), .a_0_(temp_add_fir[48]), .product_31_(
        mul_add_fir[123]), .product_30_(mul_add_fir[122]), .product_29_(
        mul_add_fir[121]), .product_28_(mul_add_fir[120]), .product_27_(
        mul_add_fir[119]), .product_26_(mul_add_fir[118]), .product_25_(
        mul_add_fir[117]), .product_24_(mul_add_fir[116]), .product_23_(
        mul_add_fir[115]), .product_22_(mul_add_fir[114]), .product_21_(
        mul_add_fir[113]), .product_20_(mul_add_fir[112]), .product_19_(
        mul_add_fir[111]), .product_18_(mul_add_fir[110]), .product_17_(
        mul_add_fir[109]), .product_16_(mul_add_fir[108]), .product_15_(
        mul_add_fir[107]), .product_14_(mul_add_fir[106]), .product_13_(
        mul_add_fir[105]), .product_12_(mul_add_fir[104]), .product_11_(
        mul_add_fir[103]), .product_10_(mul_add_fir[102]), .product_9_(
        mul_add_fir[101]), .product_8_(mul_add_fir[100]), .product_7_(
        mul_add_fir[99]), .product_6_(mul_add_fir[98]), .product_5_(
        mul_add_fir[97]), .product_4_(mul_add_fir[96]), .product_3_(
        mul_add_fir[95]), .product_2_(mul_add_fir[94]), .product_1_(
        mul_add_fir[93]) );
  FIR_FILTER2_DW_mult_uns_2 mult_126 ( .a_16_(temp_add_fir[47]), .a_14_(
        temp_add_fir[46]), .a_13_(temp_add_fir[45]), .a_12_(temp_add_fir[44]), 
        .a_11_(temp_add_fir[43]), .a_10_(temp_add_fir[42]), .a_9_(
        temp_add_fir[41]), .a_8_(temp_add_fir[40]), .a_7_(temp_add_fir[39]), 
        .a_6_(temp_add_fir[38]), .a_5_(temp_add_fir[37]), .a_4_(
        temp_add_fir[36]), .a_3_(temp_add_fir[35]), .a_2_(temp_add_fir[34]), 
        .a_1_(temp_add_fir[33]), .a_0_(temp_add_fir[32]), .product_31_(
        mul_add_fir[92]), .product_30_(mul_add_fir[91]), .product_29_(
        mul_add_fir[90]), .product_28_(mul_add_fir[89]), .product_27_(
        mul_add_fir[88]), .product_26_(mul_add_fir[87]), .product_25_(
        mul_add_fir[86]), .product_24_(mul_add_fir[85]), .product_23_(
        mul_add_fir[84]), .product_22_(mul_add_fir[83]), .product_21_(
        mul_add_fir[82]), .product_20_(mul_add_fir[81]), .product_19_(
        mul_add_fir[80]), .product_18_(mul_add_fir[79]), .product_17_(
        mul_add_fir[78]), .product_16_(mul_add_fir[77]), .product_15_(
        mul_add_fir[76]), .product_14_(mul_add_fir[75]), .product_13_(
        mul_add_fir[74]), .product_12_(mul_add_fir[73]), .product_11_(
        mul_add_fir[72]), .product_10_(mul_add_fir[71]), .product_9_(
        mul_add_fir[70]), .product_8_(mul_add_fir[69]), .product_7_(
        mul_add_fir[68]), .product_6_(mul_add_fir[67]), .product_5_(
        mul_add_fir[66]), .product_4_(mul_add_fir[65]), .product_3_(
        mul_add_fir[64]), .product_2_(mul_add_fir[63]) );
  FIR_FILTER2_DW_mult_uns_1 mult_127 ( .a_15_(temp_add_fir[31]), .a_14_(
        temp_add_fir[30]), .a_13_(temp_add_fir[29]), .a_12_(temp_add_fir[28]), 
        .a_11_(temp_add_fir[27]), .a_10_(temp_add_fir[26]), .a_9_(
        temp_add_fir[25]), .a_8_(temp_add_fir[24]), .a_7_(temp_add_fir[23]), 
        .a_6_(temp_add_fir[22]), .a_5_(temp_add_fir[21]), .a_4_(
        temp_add_fir[20]), .a_3_(temp_add_fir[19]), .a_2_(temp_add_fir[18]), 
        .a_1_(temp_add_fir[17]), .a_0_(temp_add_fir[16]), .product_31_(
        mul_add_fir[62]), .product_30_(mul_add_fir[61]), .product_29_(
        mul_add_fir[60]), .product_28_(mul_add_fir[59]), .product_27_(
        mul_add_fir[58]), .product_26_(mul_add_fir[57]), .product_25_(
        mul_add_fir[56]), .product_24_(mul_add_fir[55]), .product_23_(
        mul_add_fir[54]), .product_22_(mul_add_fir[53]), .product_21_(
        mul_add_fir[52]), .product_20_(mul_add_fir[51]), .product_19_(
        mul_add_fir[50]), .product_18_(mul_add_fir[49]), .product_17_(
        mul_add_fir[48]), .product_16_(mul_add_fir[47]), .product_15_(
        mul_add_fir[46]), .product_14_(mul_add_fir[45]), .product_13_(
        mul_add_fir[44]), .product_12_(mul_add_fir[43]), .product_11_(
        mul_add_fir[42]), .product_10_(mul_add_fir[41]), .product_9_(
        mul_add_fir[40]), .product_8_(mul_add_fir[39]), .product_7_(
        mul_add_fir[38]), .product_6_(mul_add_fir[37]), .product_5_(
        mul_add_fir[36]), .product_4_(mul_add_fir[35]), .product_3_(
        mul_add_fir[34]), .product_2_(mul_add_fir[33]), .product_1_(
        mul_add_fir[32]) );
  FIR_FILTER2_DW_mult_uns_0 mult_128 ( .a_15_(temp_add_fir[15]), .a_14_(
        temp_add_fir[14]), .a_13_(temp_add_fir[13]), .a_12_(temp_add_fir[12]), 
        .a_11_(temp_add_fir[11]), .a_10_(temp_add_fir[10]), .a_9_(
        temp_add_fir[9]), .a_8_(temp_add_fir[8]), .a_7_(temp_add_fir[7]), 
        .a_6_(temp_add_fir[6]), .a_5_(temp_add_fir[5]), .a_4_(temp_add_fir[4]), 
        .a_3_(temp_add_fir[3]), .a_2_(temp_add_fir[2]), .a_1_(temp_add_fir[1]), 
        .a_0_(temp_add_fir[0]), .product_31_(mul_add_fir[31]), .product_30_(
        mul_add_fir[30]), .product_29_(mul_add_fir[29]), .product_28_(
        mul_add_fir[28]), .product_27_(mul_add_fir[27]), .product_26_(
        mul_add_fir[26]), .product_25_(mul_add_fir[25]), .product_24_(
        mul_add_fir[24]), .product_23_(mul_add_fir[23]), .product_22_(
        mul_add_fir[22]), .product_21_(mul_add_fir[21]), .product_20_(
        mul_add_fir[20]), .product_19_(mul_add_fir[19]), .product_18_(
        mul_add_fir[18]), .product_17_(mul_add_fir[17]), .product_16_(
        mul_add_fir[16]), .product_15_(mul_add_fir[15]), .product_14_(
        mul_add_fir[14]), .product_13_(mul_add_fir[13]), .product_12_(
        mul_add_fir[12]), .product_11_(mul_add_fir[11]), .product_10_(
        mul_add_fir[10]), .product_9_(mul_add_fir[9]), .product_8_(
        mul_add_fir[8]), .product_7_(mul_add_fir[7]), .product_6_(
        mul_add_fir[6]), .product_5_(mul_add_fir[5]), .product_4_(
        mul_add_fir[4]), .product_3_(mul_add_fir[3]), .product_2_(
        mul_add_fir[2]), .product_1_(mul_add_fir[1]), .product_0_(
        mul_add_fir[0]) );
  ADDFXL mult_120_U34 ( .A(temp_add_fir[129]), .B(n750), .CI(mult_120_n29), 
        .CO(mult_120_n28), .S(mul_add_fir[252]) );
  ADDFXL mult_120_U33 ( .A(temp_add_fir[130]), .B(n760), .CI(mult_120_n28), 
        .CO(mult_120_n27), .S(mul_add_fir[253]) );
  ADDFXL mult_120_U32 ( .A(temp_add_fir[131]), .B(n770), .CI(mult_120_n27), 
        .CO(mult_120_n26), .S(mul_add_fir[254]) );
  ADDFXL mult_120_U31 ( .A(temp_add_fir[132]), .B(n780), .CI(mult_120_n26), 
        .CO(mult_120_n25), .S(mul_add_fir[255]) );
  ADDFXL mult_120_U30 ( .A(temp_add_fir[133]), .B(n790), .CI(mult_120_n25), 
        .CO(mult_120_n24), .S(mul_add_fir[256]) );
  ADDFXL mult_120_U29 ( .A(temp_add_fir[134]), .B(n800), .CI(mult_120_n24), 
        .CO(mult_120_n23), .S(mul_add_fir[257]) );
  ADDFXL mult_120_U28 ( .A(temp_add_fir[135]), .B(n810), .CI(mult_120_n23), 
        .CO(mult_120_n22), .S(mul_add_fir[258]) );
  ADDFXL mult_120_U27 ( .A(temp_add_fir[136]), .B(n820), .CI(mult_120_n22), 
        .CO(mult_120_n21), .S(mul_add_fir[259]) );
  ADDFXL mult_120_U26 ( .A(temp_add_fir[137]), .B(n830), .CI(mult_120_n21), 
        .CO(mult_120_n20), .S(mul_add_fir[260]) );
  ADDFXL mult_120_U25 ( .A(temp_add_fir[138]), .B(n840), .CI(mult_120_n20), 
        .CO(mult_120_n19), .S(mul_add_fir[261]) );
  ADDFXL mult_120_U24 ( .A(temp_add_fir[139]), .B(n850), .CI(mult_120_n19), 
        .CO(mult_120_n18), .S(mul_add_fir[262]) );
  ADDFXL mult_120_U23 ( .A(n860), .B(temp_add_fir[140]), .CI(mult_120_n18), 
        .CO(mult_120_n17), .S(mul_add_fir[263]) );
  ADDFXL mult_120_U22 ( .A(n890), .B(temp_add_fir[138]), .CI(mult_120_n17), 
        .CO(mult_120_n16), .S(mul_add_fir[264]) );
  ADDFXL mult_120_U21 ( .A(n870), .B(temp_add_fir[139]), .CI(mult_120_n16), 
        .CO(mult_120_n15), .S(mul_add_fir[265]) );
  ADDFXL mult_120_U20 ( .A(temp_add_fir[140]), .B(n880), .CI(mult_120_n15), 
        .CO(mult_120_n14), .S(mul_add_fir[266]) );
  DFFQX1 fir_data_reg_1__15_ ( .D(fir_data[511]), .CK(clk), .Q(fir_data[495])
         );
  DFFQX1 fir_data_reg_1__14_ ( .D(fir_data[510]), .CK(clk), .Q(fir_data[494])
         );
  DFFQX1 fir_data_reg_1__13_ ( .D(fir_data[509]), .CK(clk), .Q(fir_data[493])
         );
  DFFQX1 fir_data_reg_1__12_ ( .D(fir_data[508]), .CK(clk), .Q(fir_data[492])
         );
  DFFQX1 fir_data_reg_2__15_ ( .D(fir_data[495]), .CK(clk), .Q(fir_data[479])
         );
  DFFQX1 fir_data_reg_2__14_ ( .D(fir_data[494]), .CK(clk), .Q(fir_data[478])
         );
  DFFQX1 fir_data_reg_2__13_ ( .D(fir_data[493]), .CK(clk), .Q(fir_data[477])
         );
  DFFQX1 fir_data_reg_2__12_ ( .D(fir_data[492]), .CK(clk), .Q(fir_data[476])
         );
  DFFQX1 fir_data_reg_3__15_ ( .D(fir_data[479]), .CK(clk), .Q(fir_data[463])
         );
  DFFQX1 fir_data_reg_3__14_ ( .D(fir_data[478]), .CK(clk), .Q(fir_data[462])
         );
  DFFQX1 fir_data_reg_3__13_ ( .D(fir_data[477]), .CK(clk), .Q(fir_data[461])
         );
  DFFQX1 fir_data_reg_3__12_ ( .D(fir_data[476]), .CK(clk), .Q(fir_data[460])
         );
  DFFQX1 fir_data_reg_4__15_ ( .D(fir_data[463]), .CK(clk), .Q(fir_data[447])
         );
  DFFQX1 fir_data_reg_4__14_ ( .D(fir_data[462]), .CK(clk), .Q(fir_data[446])
         );
  DFFQX1 fir_data_reg_4__13_ ( .D(fir_data[461]), .CK(clk), .Q(fir_data[445])
         );
  DFFQX1 fir_data_reg_4__12_ ( .D(fir_data[460]), .CK(clk), .Q(fir_data[444])
         );
  DFFQX1 fir_data_reg_5__15_ ( .D(fir_data[447]), .CK(clk), .Q(fir_data[431])
         );
  DFFQX1 fir_data_reg_5__14_ ( .D(fir_data[446]), .CK(clk), .Q(fir_data[430])
         );
  DFFQX1 fir_data_reg_5__13_ ( .D(fir_data[445]), .CK(clk), .Q(fir_data[429])
         );
  DFFQX1 fir_data_reg_5__12_ ( .D(fir_data[444]), .CK(clk), .Q(fir_data[428])
         );
  DFFQX1 fir_data_reg_6__15_ ( .D(fir_data[431]), .CK(clk), .Q(fir_data[415])
         );
  DFFQX1 fir_data_reg_6__14_ ( .D(fir_data[430]), .CK(clk), .Q(fir_data[414])
         );
  DFFQX1 fir_data_reg_6__13_ ( .D(fir_data[429]), .CK(clk), .Q(fir_data[413])
         );
  DFFQX1 fir_data_reg_6__12_ ( .D(fir_data[428]), .CK(clk), .Q(fir_data[412])
         );
  DFFQX1 fir_data_reg_7__15_ ( .D(fir_data[415]), .CK(clk), .Q(fir_data[399])
         );
  DFFQX1 fir_data_reg_7__14_ ( .D(fir_data[414]), .CK(clk), .Q(fir_data[398])
         );
  DFFQX1 fir_data_reg_7__13_ ( .D(fir_data[413]), .CK(clk), .Q(fir_data[397])
         );
  DFFQX1 fir_data_reg_7__12_ ( .D(fir_data[412]), .CK(clk), .Q(fir_data[396])
         );
  DFFQX1 fir_data_reg_8__15_ ( .D(fir_data[399]), .CK(clk), .Q(fir_data[383])
         );
  DFFQX1 fir_data_reg_8__14_ ( .D(fir_data[398]), .CK(clk), .Q(fir_data[382])
         );
  DFFQX1 fir_data_reg_8__13_ ( .D(fir_data[397]), .CK(clk), .Q(fir_data[381])
         );
  DFFQX1 fir_data_reg_8__12_ ( .D(fir_data[396]), .CK(clk), .Q(fir_data[380])
         );
  DFFQX1 fir_data_reg_9__15_ ( .D(fir_data[383]), .CK(clk), .Q(fir_data[367])
         );
  DFFQX1 fir_data_reg_9__14_ ( .D(fir_data[382]), .CK(clk), .Q(fir_data[366])
         );
  DFFQX1 fir_data_reg_9__13_ ( .D(fir_data[381]), .CK(clk), .Q(fir_data[365])
         );
  DFFQX1 fir_data_reg_9__12_ ( .D(fir_data[380]), .CK(clk), .Q(fir_data[364])
         );
  DFFQX1 fir_data_reg_10__15_ ( .D(fir_data[367]), .CK(clk), .Q(fir_data[351])
         );
  DFFQX1 fir_data_reg_10__14_ ( .D(fir_data[366]), .CK(clk), .Q(fir_data[350])
         );
  DFFQX1 fir_data_reg_10__13_ ( .D(fir_data[365]), .CK(clk), .Q(fir_data[349])
         );
  DFFQX1 fir_data_reg_10__12_ ( .D(fir_data[364]), .CK(clk), .Q(fir_data[348])
         );
  DFFQX1 fir_data_reg_11__15_ ( .D(fir_data[351]), .CK(clk), .Q(fir_data[335])
         );
  DFFQX1 fir_data_reg_11__14_ ( .D(fir_data[350]), .CK(clk), .Q(fir_data[334])
         );
  DFFQX1 fir_data_reg_11__13_ ( .D(fir_data[349]), .CK(clk), .Q(fir_data[333])
         );
  DFFQX1 fir_data_reg_11__12_ ( .D(fir_data[348]), .CK(clk), .Q(fir_data[332])
         );
  DFFQX1 fir_data_reg_12__15_ ( .D(fir_data[335]), .CK(clk), .Q(fir_data[319])
         );
  DFFQX1 fir_data_reg_12__14_ ( .D(fir_data[334]), .CK(clk), .Q(fir_data[318])
         );
  DFFQX1 fir_data_reg_12__13_ ( .D(fir_data[333]), .CK(clk), .Q(fir_data[317])
         );
  DFFQX1 fir_data_reg_12__12_ ( .D(fir_data[332]), .CK(clk), .Q(fir_data[316])
         );
  DFFQX1 fir_data_reg_13__15_ ( .D(fir_data[319]), .CK(clk), .Q(fir_data[303])
         );
  DFFQX1 fir_data_reg_13__14_ ( .D(fir_data[318]), .CK(clk), .Q(fir_data[302])
         );
  DFFQX1 fir_data_reg_13__13_ ( .D(fir_data[317]), .CK(clk), .Q(fir_data[301])
         );
  DFFQX1 fir_data_reg_13__12_ ( .D(fir_data[316]), .CK(clk), .Q(fir_data[300])
         );
  DFFQX1 fir_data_reg_14__15_ ( .D(fir_data[303]), .CK(clk), .Q(fir_data[287])
         );
  DFFQX1 fir_data_reg_14__14_ ( .D(fir_data[302]), .CK(clk), .Q(fir_data[286])
         );
  DFFQX1 fir_data_reg_14__13_ ( .D(fir_data[301]), .CK(clk), .Q(fir_data[285])
         );
  DFFQX1 fir_data_reg_14__12_ ( .D(fir_data[300]), .CK(clk), .Q(fir_data[284])
         );
  DFFQX1 fir_data_reg_15__15_ ( .D(fir_data[287]), .CK(clk), .Q(fir_data[271])
         );
  DFFQX1 fir_data_reg_15__14_ ( .D(fir_data[286]), .CK(clk), .Q(fir_data[270])
         );
  DFFQX1 fir_data_reg_15__13_ ( .D(fir_data[285]), .CK(clk), .Q(fir_data[269])
         );
  DFFQX1 fir_data_reg_15__12_ ( .D(fir_data[284]), .CK(clk), .Q(fir_data[268])
         );
  DFFTRX1 fir_data_reg_0__15_ ( .D(data[15]), .RN(n56), .CK(clk), .Q(
        fir_data[511]) );
  DFFTRX1 fir_data_reg_0__14_ ( .D(data[14]), .RN(n56), .CK(clk), .Q(
        fir_data[510]) );
  DFFTRX1 fir_data_reg_0__13_ ( .D(data[13]), .RN(n56), .CK(clk), .Q(
        fir_data[509]) );
  DFFQX1 fir_data_reg_31__15_ ( .D(fir_data[31]), .CK(clk), .Q(fir_data[15])
         );
  DFFQX1 fir_data_reg_31__14_ ( .D(fir_data[30]), .CK(clk), .Q(fir_data[14])
         );
  DFFQX1 fir_data_reg_31__13_ ( .D(fir_data[29]), .CK(clk), .Q(fir_data[13])
         );
  DFFQX1 fir_data_reg_31__12_ ( .D(fir_data[28]), .CK(clk), .Q(fir_data[12])
         );
  DFFQX1 fir_data_reg_16__15_ ( .D(fir_data[271]), .CK(clk), .Q(fir_data[255])
         );
  DFFQX1 fir_data_reg_16__14_ ( .D(fir_data[270]), .CK(clk), .Q(fir_data[254])
         );
  DFFQX1 fir_data_reg_16__13_ ( .D(fir_data[269]), .CK(clk), .Q(fir_data[253])
         );
  DFFQX1 fir_data_reg_16__12_ ( .D(fir_data[268]), .CK(clk), .Q(fir_data[252])
         );
  DFFQX1 fir_data_reg_17__15_ ( .D(fir_data[255]), .CK(clk), .Q(fir_data[239])
         );
  DFFQX1 fir_data_reg_17__14_ ( .D(fir_data[254]), .CK(clk), .Q(fir_data[238])
         );
  DFFQX1 fir_data_reg_17__13_ ( .D(fir_data[253]), .CK(clk), .Q(fir_data[237])
         );
  DFFQX1 fir_data_reg_17__12_ ( .D(fir_data[252]), .CK(clk), .Q(fir_data[236])
         );
  DFFQX1 fir_data_reg_18__15_ ( .D(fir_data[239]), .CK(clk), .Q(fir_data[223])
         );
  DFFQX1 fir_data_reg_18__14_ ( .D(fir_data[238]), .CK(clk), .Q(fir_data[222])
         );
  DFFQX1 fir_data_reg_18__13_ ( .D(fir_data[237]), .CK(clk), .Q(fir_data[221])
         );
  DFFQX1 fir_data_reg_18__12_ ( .D(fir_data[236]), .CK(clk), .Q(fir_data[220])
         );
  DFFQX1 fir_data_reg_19__15_ ( .D(fir_data[223]), .CK(clk), .Q(fir_data[207])
         );
  DFFQX1 fir_data_reg_19__14_ ( .D(fir_data[222]), .CK(clk), .Q(fir_data[206])
         );
  DFFQX1 fir_data_reg_19__13_ ( .D(fir_data[221]), .CK(clk), .Q(fir_data[205])
         );
  DFFQX1 fir_data_reg_19__12_ ( .D(fir_data[220]), .CK(clk), .Q(fir_data[204])
         );
  DFFQX1 fir_data_reg_20__15_ ( .D(fir_data[207]), .CK(clk), .Q(fir_data[191])
         );
  DFFQX1 fir_data_reg_20__14_ ( .D(fir_data[206]), .CK(clk), .Q(fir_data[190])
         );
  DFFQX1 fir_data_reg_20__13_ ( .D(fir_data[205]), .CK(clk), .Q(fir_data[189])
         );
  DFFQX1 fir_data_reg_20__12_ ( .D(fir_data[204]), .CK(clk), .Q(fir_data[188])
         );
  DFFQX1 fir_data_reg_21__15_ ( .D(fir_data[191]), .CK(clk), .Q(fir_data[175])
         );
  DFFQX1 fir_data_reg_21__14_ ( .D(fir_data[190]), .CK(clk), .Q(fir_data[174])
         );
  DFFQX1 fir_data_reg_21__13_ ( .D(fir_data[189]), .CK(clk), .Q(fir_data[173])
         );
  DFFQX1 fir_data_reg_21__12_ ( .D(fir_data[188]), .CK(clk), .Q(fir_data[172])
         );
  DFFQX1 fir_data_reg_22__15_ ( .D(fir_data[175]), .CK(clk), .Q(fir_data[159])
         );
  DFFQX1 fir_data_reg_22__14_ ( .D(fir_data[174]), .CK(clk), .Q(fir_data[158])
         );
  DFFQX1 fir_data_reg_22__13_ ( .D(fir_data[173]), .CK(clk), .Q(fir_data[157])
         );
  DFFQX1 fir_data_reg_22__12_ ( .D(fir_data[172]), .CK(clk), .Q(fir_data[156])
         );
  DFFQX1 fir_data_reg_23__15_ ( .D(fir_data[159]), .CK(clk), .Q(fir_data[143])
         );
  DFFQX1 fir_data_reg_23__14_ ( .D(fir_data[158]), .CK(clk), .Q(fir_data[142])
         );
  DFFQX1 fir_data_reg_23__13_ ( .D(fir_data[157]), .CK(clk), .Q(fir_data[141])
         );
  DFFQX1 fir_data_reg_23__12_ ( .D(fir_data[156]), .CK(clk), .Q(fir_data[140])
         );
  DFFQX1 fir_data_reg_24__15_ ( .D(fir_data[143]), .CK(clk), .Q(fir_data[127])
         );
  DFFQX1 fir_data_reg_24__14_ ( .D(fir_data[142]), .CK(clk), .Q(fir_data[126])
         );
  DFFQX1 fir_data_reg_24__13_ ( .D(fir_data[141]), .CK(clk), .Q(fir_data[125])
         );
  DFFQX1 fir_data_reg_24__12_ ( .D(fir_data[140]), .CK(clk), .Q(fir_data[124])
         );
  DFFQX1 fir_data_reg_25__15_ ( .D(fir_data[127]), .CK(clk), .Q(fir_data[111])
         );
  DFFQX1 fir_data_reg_25__14_ ( .D(fir_data[126]), .CK(clk), .Q(fir_data[110])
         );
  DFFQX1 fir_data_reg_25__13_ ( .D(fir_data[125]), .CK(clk), .Q(fir_data[109])
         );
  DFFQX1 fir_data_reg_25__12_ ( .D(fir_data[124]), .CK(clk), .Q(fir_data[108])
         );
  DFFQX1 fir_data_reg_26__15_ ( .D(fir_data[111]), .CK(clk), .Q(fir_data[95])
         );
  DFFQX1 fir_data_reg_26__14_ ( .D(fir_data[110]), .CK(clk), .Q(fir_data[94])
         );
  DFFQX1 fir_data_reg_26__13_ ( .D(fir_data[109]), .CK(clk), .Q(fir_data[93])
         );
  DFFQX1 fir_data_reg_26__12_ ( .D(fir_data[108]), .CK(clk), .Q(fir_data[92])
         );
  DFFQX1 fir_data_reg_27__15_ ( .D(fir_data[95]), .CK(clk), .Q(fir_data[79])
         );
  DFFQX1 fir_data_reg_27__14_ ( .D(fir_data[94]), .CK(clk), .Q(fir_data[78])
         );
  DFFQX1 fir_data_reg_27__13_ ( .D(fir_data[93]), .CK(clk), .Q(fir_data[77])
         );
  DFFQX1 fir_data_reg_27__12_ ( .D(fir_data[92]), .CK(clk), .Q(fir_data[76])
         );
  DFFQX1 fir_data_reg_28__15_ ( .D(fir_data[79]), .CK(clk), .Q(fir_data[63])
         );
  DFFQX1 fir_data_reg_28__14_ ( .D(fir_data[78]), .CK(clk), .Q(fir_data[62])
         );
  DFFQX1 fir_data_reg_28__13_ ( .D(fir_data[77]), .CK(clk), .Q(fir_data[61])
         );
  DFFQX1 fir_data_reg_28__12_ ( .D(fir_data[76]), .CK(clk), .Q(fir_data[60])
         );
  DFFQX1 fir_data_reg_29__15_ ( .D(fir_data[63]), .CK(clk), .Q(fir_data[47])
         );
  DFFQX1 fir_data_reg_29__14_ ( .D(fir_data[62]), .CK(clk), .Q(fir_data[46])
         );
  DFFQX1 fir_data_reg_29__13_ ( .D(fir_data[61]), .CK(clk), .Q(fir_data[45])
         );
  DFFQX1 fir_data_reg_29__12_ ( .D(fir_data[60]), .CK(clk), .Q(fir_data[44])
         );
  DFFQX1 fir_data_reg_30__15_ ( .D(fir_data[47]), .CK(clk), .Q(fir_data[31])
         );
  DFFQX1 fir_data_reg_30__14_ ( .D(fir_data[46]), .CK(clk), .Q(fir_data[30])
         );
  DFFQX1 fir_data_reg_30__13_ ( .D(fir_data[45]), .CK(clk), .Q(fir_data[29])
         );
  DFFQX1 fir_data_reg_30__12_ ( .D(fir_data[44]), .CK(clk), .Q(fir_data[28])
         );
  DFFQX1 temp_mul_add_fir_reg_0__31_ ( .D(mul_add_fir[487]), .CK(clk), .Q(
        temp_mul_add_fir[511]) );
  DFFQX1 temp_mul_add_fir_reg_0__30_ ( .D(mul_add_fir[486]), .CK(clk), .Q(
        temp_mul_add_fir[510]) );
  DFFQX1 temp_mul_add_fir_reg_0__29_ ( .D(mul_add_fir[485]), .CK(clk), .Q(
        temp_mul_add_fir[509]) );
  DFFQX1 temp_mul_add_fir_reg_0__28_ ( .D(mul_add_fir[484]), .CK(clk), .Q(
        temp_mul_add_fir[508]) );
  DFFQX1 temp_mul_add_fir_reg_2__31_ ( .D(mul_add_fir[425]), .CK(clk), .Q(
        temp_mul_add_fir[447]) );
  DFFQX1 temp_mul_add_fir_reg_2__30_ ( .D(mul_add_fir[424]), .CK(clk), .Q(
        temp_mul_add_fir[446]) );
  DFFQX1 temp_mul_add_fir_reg_2__29_ ( .D(mul_add_fir[423]), .CK(clk), .Q(
        temp_mul_add_fir[445]) );
  DFFQX1 temp_mul_add_fir_reg_2__28_ ( .D(mul_add_fir[422]), .CK(clk), .Q(
        temp_mul_add_fir[444]) );
  DFFQX1 temp_mul_add_fir_reg_4__31_ ( .D(mul_add_fir[361]), .CK(clk), .Q(
        temp_mul_add_fir[383]) );
  DFFQX1 temp_mul_add_fir_reg_4__30_ ( .D(mul_add_fir[360]), .CK(clk), .Q(
        temp_mul_add_fir[382]) );
  DFFQX1 temp_mul_add_fir_reg_4__29_ ( .D(mul_add_fir[359]), .CK(clk), .Q(
        temp_mul_add_fir[381]) );
  DFFQX1 temp_mul_add_fir_reg_4__28_ ( .D(mul_add_fir[358]), .CK(clk), .Q(
        temp_mul_add_fir[380]) );
  DFFQX1 temp_mul_add_fir_reg_6__31_ ( .D(mul_add_fir[298]), .CK(clk), .Q(
        temp_mul_add_fir[319]) );
  DFFQX1 temp_mul_add_fir_reg_6__30_ ( .D(mul_add_fir[297]), .CK(clk), .Q(
        temp_mul_add_fir[318]) );
  DFFQX1 temp_mul_add_fir_reg_6__29_ ( .D(mul_add_fir[296]), .CK(clk), .Q(
        temp_mul_add_fir[317]) );
  DFFQX1 temp_mul_add_fir_reg_6__28_ ( .D(mul_add_fir[295]), .CK(clk), .Q(
        temp_mul_add_fir[316]) );
  DFFQX1 temp_mul_add_fir_reg_8__31_ ( .D(mul_add_fir[247]), .CK(clk), .Q(
        temp_mul_add_fir[255]) );
  DFFQX1 temp_mul_add_fir_reg_8__30_ ( .D(mul_add_fir[246]), .CK(clk), .Q(
        temp_mul_add_fir[254]) );
  DFFQX1 temp_mul_add_fir_reg_8__29_ ( .D(mul_add_fir[245]), .CK(clk), .Q(
        temp_mul_add_fir[253]) );
  DFFQX1 temp_mul_add_fir_reg_8__28_ ( .D(mul_add_fir[244]), .CK(clk), .Q(
        temp_mul_add_fir[252]) );
  DFFQX1 temp_mul_add_fir_reg_10__31_ ( .D(mul_add_fir[184]), .CK(clk), .Q(
        temp_mul_add_fir[191]) );
  DFFQX1 temp_mul_add_fir_reg_10__30_ ( .D(mul_add_fir[183]), .CK(clk), .Q(
        temp_mul_add_fir[190]) );
  DFFQX1 temp_mul_add_fir_reg_10__29_ ( .D(mul_add_fir[182]), .CK(clk), .Q(
        temp_mul_add_fir[189]) );
  DFFQX1 temp_mul_add_fir_reg_10__28_ ( .D(mul_add_fir[181]), .CK(clk), .Q(
        temp_mul_add_fir[188]) );
  DFFQX1 temp_mul_add_fir_reg_12__31_ ( .D(mul_add_fir[123]), .CK(clk), .Q(
        temp_mul_add_fir[127]) );
  DFFQX1 temp_mul_add_fir_reg_12__30_ ( .D(mul_add_fir[122]), .CK(clk), .Q(
        temp_mul_add_fir[126]) );
  DFFQX1 temp_mul_add_fir_reg_12__29_ ( .D(mul_add_fir[121]), .CK(clk), .Q(
        temp_mul_add_fir[125]) );
  DFFQX1 temp_mul_add_fir_reg_12__28_ ( .D(mul_add_fir[120]), .CK(clk), .Q(
        temp_mul_add_fir[124]) );
  DFFQX1 temp_mul_add_fir_reg_14__31_ ( .D(mul_add_fir[62]), .CK(clk), .Q(
        temp_mul_add_fir[63]) );
  DFFQX1 temp_mul_add_fir_reg_14__30_ ( .D(mul_add_fir[61]), .CK(clk), .Q(
        temp_mul_add_fir[62]) );
  DFFQX1 temp_mul_add_fir_reg_14__29_ ( .D(mul_add_fir[60]), .CK(clk), .Q(
        temp_mul_add_fir[61]) );
  DFFQX1 temp_mul_add_fir_reg_14__28_ ( .D(mul_add_fir[59]), .CK(clk), .Q(
        temp_mul_add_fir[60]) );
  DFFQX1 fir_data_reg_1__11_ ( .D(fir_data[507]), .CK(clk), .Q(fir_data[491])
         );
  DFFQX1 fir_data_reg_1__10_ ( .D(fir_data[506]), .CK(clk), .Q(fir_data[490])
         );
  DFFQX1 fir_data_reg_1__9_ ( .D(fir_data[505]), .CK(clk), .Q(fir_data[489])
         );
  DFFQX1 fir_data_reg_1__8_ ( .D(fir_data[504]), .CK(clk), .Q(fir_data[488])
         );
  DFFQX1 fir_data_reg_1__7_ ( .D(fir_data[503]), .CK(clk), .Q(fir_data[487])
         );
  DFFQX1 fir_data_reg_1__6_ ( .D(fir_data[502]), .CK(clk), .Q(fir_data[486])
         );
  DFFQX1 fir_data_reg_1__5_ ( .D(fir_data[501]), .CK(clk), .Q(fir_data[485])
         );
  DFFQX1 fir_data_reg_1__4_ ( .D(fir_data[500]), .CK(clk), .Q(fir_data[484])
         );
  DFFQX1 fir_data_reg_2__11_ ( .D(fir_data[491]), .CK(clk), .Q(fir_data[475])
         );
  DFFQX1 fir_data_reg_2__10_ ( .D(fir_data[490]), .CK(clk), .Q(fir_data[474])
         );
  DFFQX1 fir_data_reg_2__9_ ( .D(fir_data[489]), .CK(clk), .Q(fir_data[473])
         );
  DFFQX1 fir_data_reg_2__8_ ( .D(fir_data[488]), .CK(clk), .Q(fir_data[472])
         );
  DFFQX1 fir_data_reg_2__7_ ( .D(fir_data[487]), .CK(clk), .Q(fir_data[471])
         );
  DFFQX1 fir_data_reg_2__6_ ( .D(fir_data[486]), .CK(clk), .Q(fir_data[470])
         );
  DFFQX1 fir_data_reg_2__5_ ( .D(fir_data[485]), .CK(clk), .Q(fir_data[469])
         );
  DFFQX1 fir_data_reg_2__4_ ( .D(fir_data[484]), .CK(clk), .Q(fir_data[468])
         );
  DFFQX1 fir_data_reg_3__11_ ( .D(fir_data[475]), .CK(clk), .Q(fir_data[459])
         );
  DFFQX1 fir_data_reg_3__10_ ( .D(fir_data[474]), .CK(clk), .Q(fir_data[458])
         );
  DFFQX1 fir_data_reg_3__9_ ( .D(fir_data[473]), .CK(clk), .Q(fir_data[457])
         );
  DFFQX1 fir_data_reg_3__8_ ( .D(fir_data[472]), .CK(clk), .Q(fir_data[456])
         );
  DFFQX1 fir_data_reg_3__7_ ( .D(fir_data[471]), .CK(clk), .Q(fir_data[455])
         );
  DFFQX1 fir_data_reg_3__6_ ( .D(fir_data[470]), .CK(clk), .Q(fir_data[454])
         );
  DFFQX1 fir_data_reg_3__5_ ( .D(fir_data[469]), .CK(clk), .Q(fir_data[453])
         );
  DFFQX1 fir_data_reg_3__4_ ( .D(fir_data[468]), .CK(clk), .Q(fir_data[452])
         );
  DFFQX1 fir_data_reg_4__11_ ( .D(fir_data[459]), .CK(clk), .Q(fir_data[443])
         );
  DFFQX1 fir_data_reg_4__10_ ( .D(fir_data[458]), .CK(clk), .Q(fir_data[442])
         );
  DFFQX1 fir_data_reg_4__9_ ( .D(fir_data[457]), .CK(clk), .Q(fir_data[441])
         );
  DFFQX1 fir_data_reg_4__8_ ( .D(fir_data[456]), .CK(clk), .Q(fir_data[440])
         );
  DFFQX1 fir_data_reg_4__7_ ( .D(fir_data[455]), .CK(clk), .Q(fir_data[439])
         );
  DFFQX1 fir_data_reg_4__6_ ( .D(fir_data[454]), .CK(clk), .Q(fir_data[438])
         );
  DFFQX1 fir_data_reg_4__5_ ( .D(fir_data[453]), .CK(clk), .Q(fir_data[437])
         );
  DFFQX1 fir_data_reg_4__4_ ( .D(fir_data[452]), .CK(clk), .Q(fir_data[436])
         );
  DFFQX1 fir_data_reg_5__11_ ( .D(fir_data[443]), .CK(clk), .Q(fir_data[427])
         );
  DFFQX1 fir_data_reg_5__10_ ( .D(fir_data[442]), .CK(clk), .Q(fir_data[426])
         );
  DFFQX1 fir_data_reg_5__9_ ( .D(fir_data[441]), .CK(clk), .Q(fir_data[425])
         );
  DFFQX1 fir_data_reg_5__8_ ( .D(fir_data[440]), .CK(clk), .Q(fir_data[424])
         );
  DFFQX1 fir_data_reg_5__7_ ( .D(fir_data[439]), .CK(clk), .Q(fir_data[423])
         );
  DFFQX1 fir_data_reg_5__6_ ( .D(fir_data[438]), .CK(clk), .Q(fir_data[422])
         );
  DFFQX1 fir_data_reg_5__5_ ( .D(fir_data[437]), .CK(clk), .Q(fir_data[421])
         );
  DFFQX1 fir_data_reg_5__4_ ( .D(fir_data[436]), .CK(clk), .Q(fir_data[420])
         );
  DFFQX1 fir_data_reg_6__11_ ( .D(fir_data[427]), .CK(clk), .Q(fir_data[411])
         );
  DFFQX1 fir_data_reg_6__10_ ( .D(fir_data[426]), .CK(clk), .Q(fir_data[410])
         );
  DFFQX1 fir_data_reg_6__9_ ( .D(fir_data[425]), .CK(clk), .Q(fir_data[409])
         );
  DFFQX1 fir_data_reg_6__8_ ( .D(fir_data[424]), .CK(clk), .Q(fir_data[408])
         );
  DFFQX1 fir_data_reg_6__7_ ( .D(fir_data[423]), .CK(clk), .Q(fir_data[407])
         );
  DFFQX1 fir_data_reg_6__6_ ( .D(fir_data[422]), .CK(clk), .Q(fir_data[406])
         );
  DFFQX1 fir_data_reg_6__5_ ( .D(fir_data[421]), .CK(clk), .Q(fir_data[405])
         );
  DFFQX1 fir_data_reg_6__4_ ( .D(fir_data[420]), .CK(clk), .Q(fir_data[404])
         );
  DFFQX1 fir_data_reg_7__11_ ( .D(fir_data[411]), .CK(clk), .Q(fir_data[395])
         );
  DFFQX1 fir_data_reg_7__10_ ( .D(fir_data[410]), .CK(clk), .Q(fir_data[394])
         );
  DFFQX1 fir_data_reg_7__9_ ( .D(fir_data[409]), .CK(clk), .Q(fir_data[393])
         );
  DFFQX1 fir_data_reg_7__8_ ( .D(fir_data[408]), .CK(clk), .Q(fir_data[392])
         );
  DFFQX1 fir_data_reg_7__7_ ( .D(fir_data[407]), .CK(clk), .Q(fir_data[391])
         );
  DFFQX1 fir_data_reg_7__6_ ( .D(fir_data[406]), .CK(clk), .Q(fir_data[390])
         );
  DFFQX1 fir_data_reg_7__5_ ( .D(fir_data[405]), .CK(clk), .Q(fir_data[389])
         );
  DFFQX1 fir_data_reg_7__4_ ( .D(fir_data[404]), .CK(clk), .Q(fir_data[388])
         );
  DFFQX1 fir_data_reg_8__11_ ( .D(fir_data[395]), .CK(clk), .Q(fir_data[379])
         );
  DFFQX1 fir_data_reg_8__10_ ( .D(fir_data[394]), .CK(clk), .Q(fir_data[378])
         );
  DFFQX1 fir_data_reg_8__9_ ( .D(fir_data[393]), .CK(clk), .Q(fir_data[377])
         );
  DFFQX1 fir_data_reg_8__8_ ( .D(fir_data[392]), .CK(clk), .Q(fir_data[376])
         );
  DFFQX1 fir_data_reg_8__7_ ( .D(fir_data[391]), .CK(clk), .Q(fir_data[375])
         );
  DFFQX1 fir_data_reg_8__6_ ( .D(fir_data[390]), .CK(clk), .Q(fir_data[374])
         );
  DFFQX1 fir_data_reg_8__5_ ( .D(fir_data[389]), .CK(clk), .Q(fir_data[373])
         );
  DFFQX1 fir_data_reg_8__4_ ( .D(fir_data[388]), .CK(clk), .Q(fir_data[372])
         );
  DFFQX1 fir_data_reg_9__11_ ( .D(fir_data[379]), .CK(clk), .Q(fir_data[363])
         );
  DFFQX1 fir_data_reg_9__10_ ( .D(fir_data[378]), .CK(clk), .Q(fir_data[362])
         );
  DFFQX1 fir_data_reg_9__9_ ( .D(fir_data[377]), .CK(clk), .Q(fir_data[361])
         );
  DFFQX1 fir_data_reg_9__8_ ( .D(fir_data[376]), .CK(clk), .Q(fir_data[360])
         );
  DFFQX1 fir_data_reg_9__7_ ( .D(fir_data[375]), .CK(clk), .Q(fir_data[359])
         );
  DFFQX1 fir_data_reg_9__6_ ( .D(fir_data[374]), .CK(clk), .Q(fir_data[358])
         );
  DFFQX1 fir_data_reg_9__5_ ( .D(fir_data[373]), .CK(clk), .Q(fir_data[357])
         );
  DFFQX1 fir_data_reg_9__4_ ( .D(fir_data[372]), .CK(clk), .Q(fir_data[356])
         );
  DFFQX1 fir_data_reg_10__11_ ( .D(fir_data[363]), .CK(clk), .Q(fir_data[347])
         );
  DFFQX1 fir_data_reg_10__10_ ( .D(fir_data[362]), .CK(clk), .Q(fir_data[346])
         );
  DFFQX1 fir_data_reg_10__9_ ( .D(fir_data[361]), .CK(clk), .Q(fir_data[345])
         );
  DFFQX1 fir_data_reg_10__8_ ( .D(fir_data[360]), .CK(clk), .Q(fir_data[344])
         );
  DFFQX1 fir_data_reg_10__7_ ( .D(fir_data[359]), .CK(clk), .Q(fir_data[343])
         );
  DFFQX1 fir_data_reg_10__6_ ( .D(fir_data[358]), .CK(clk), .Q(fir_data[342])
         );
  DFFQX1 fir_data_reg_10__5_ ( .D(fir_data[357]), .CK(clk), .Q(fir_data[341])
         );
  DFFQX1 fir_data_reg_10__4_ ( .D(fir_data[356]), .CK(clk), .Q(fir_data[340])
         );
  DFFQX1 fir_data_reg_11__11_ ( .D(fir_data[347]), .CK(clk), .Q(fir_data[331])
         );
  DFFQX1 fir_data_reg_11__10_ ( .D(fir_data[346]), .CK(clk), .Q(fir_data[330])
         );
  DFFQX1 fir_data_reg_11__9_ ( .D(fir_data[345]), .CK(clk), .Q(fir_data[329])
         );
  DFFQX1 fir_data_reg_11__8_ ( .D(fir_data[344]), .CK(clk), .Q(fir_data[328])
         );
  DFFQX1 fir_data_reg_11__7_ ( .D(fir_data[343]), .CK(clk), .Q(fir_data[327])
         );
  DFFQX1 fir_data_reg_11__6_ ( .D(fir_data[342]), .CK(clk), .Q(fir_data[326])
         );
  DFFQX1 fir_data_reg_11__5_ ( .D(fir_data[341]), .CK(clk), .Q(fir_data[325])
         );
  DFFQX1 fir_data_reg_11__4_ ( .D(fir_data[340]), .CK(clk), .Q(fir_data[324])
         );
  DFFQX1 fir_data_reg_12__11_ ( .D(fir_data[331]), .CK(clk), .Q(fir_data[315])
         );
  DFFQX1 fir_data_reg_12__10_ ( .D(fir_data[330]), .CK(clk), .Q(fir_data[314])
         );
  DFFQX1 fir_data_reg_12__9_ ( .D(fir_data[329]), .CK(clk), .Q(fir_data[313])
         );
  DFFQX1 fir_data_reg_12__8_ ( .D(fir_data[328]), .CK(clk), .Q(fir_data[312])
         );
  DFFQX1 fir_data_reg_12__7_ ( .D(fir_data[327]), .CK(clk), .Q(fir_data[311])
         );
  DFFQX1 fir_data_reg_12__6_ ( .D(fir_data[326]), .CK(clk), .Q(fir_data[310])
         );
  DFFQX1 fir_data_reg_12__5_ ( .D(fir_data[325]), .CK(clk), .Q(fir_data[309])
         );
  DFFQX1 fir_data_reg_12__4_ ( .D(fir_data[324]), .CK(clk), .Q(fir_data[308])
         );
  DFFQX1 fir_data_reg_13__11_ ( .D(fir_data[315]), .CK(clk), .Q(fir_data[299])
         );
  DFFQX1 fir_data_reg_13__10_ ( .D(fir_data[314]), .CK(clk), .Q(fir_data[298])
         );
  DFFQX1 fir_data_reg_13__9_ ( .D(fir_data[313]), .CK(clk), .Q(fir_data[297])
         );
  DFFQX1 fir_data_reg_13__8_ ( .D(fir_data[312]), .CK(clk), .Q(fir_data[296])
         );
  DFFQX1 fir_data_reg_13__7_ ( .D(fir_data[311]), .CK(clk), .Q(fir_data[295])
         );
  DFFQX1 fir_data_reg_13__6_ ( .D(fir_data[310]), .CK(clk), .Q(fir_data[294])
         );
  DFFQX1 fir_data_reg_13__5_ ( .D(fir_data[309]), .CK(clk), .Q(fir_data[293])
         );
  DFFQX1 fir_data_reg_13__4_ ( .D(fir_data[308]), .CK(clk), .Q(fir_data[292])
         );
  DFFQX1 fir_data_reg_14__11_ ( .D(fir_data[299]), .CK(clk), .Q(fir_data[283])
         );
  DFFQX1 fir_data_reg_14__10_ ( .D(fir_data[298]), .CK(clk), .Q(fir_data[282])
         );
  DFFQX1 fir_data_reg_14__9_ ( .D(fir_data[297]), .CK(clk), .Q(fir_data[281])
         );
  DFFQX1 fir_data_reg_14__8_ ( .D(fir_data[296]), .CK(clk), .Q(fir_data[280])
         );
  DFFQX1 fir_data_reg_14__7_ ( .D(fir_data[295]), .CK(clk), .Q(fir_data[279])
         );
  DFFQX1 fir_data_reg_14__6_ ( .D(fir_data[294]), .CK(clk), .Q(fir_data[278])
         );
  DFFQX1 fir_data_reg_14__5_ ( .D(fir_data[293]), .CK(clk), .Q(fir_data[277])
         );
  DFFQX1 fir_data_reg_14__4_ ( .D(fir_data[292]), .CK(clk), .Q(fir_data[276])
         );
  DFFQX1 fir_data_reg_15__11_ ( .D(fir_data[283]), .CK(clk), .Q(fir_data[267])
         );
  DFFQX1 fir_data_reg_15__10_ ( .D(fir_data[282]), .CK(clk), .Q(fir_data[266])
         );
  DFFQX1 fir_data_reg_15__9_ ( .D(fir_data[281]), .CK(clk), .Q(fir_data[265])
         );
  DFFQX1 fir_data_reg_15__8_ ( .D(fir_data[280]), .CK(clk), .Q(fir_data[264])
         );
  DFFQX1 fir_data_reg_15__7_ ( .D(fir_data[279]), .CK(clk), .Q(fir_data[263])
         );
  DFFQX1 fir_data_reg_15__6_ ( .D(fir_data[278]), .CK(clk), .Q(fir_data[262])
         );
  DFFQX1 fir_data_reg_15__5_ ( .D(fir_data[277]), .CK(clk), .Q(fir_data[261])
         );
  DFFQX1 fir_data_reg_15__4_ ( .D(fir_data[276]), .CK(clk), .Q(fir_data[260])
         );
  DFFTRX1 fir_data_reg_0__12_ ( .D(data[12]), .RN(n56), .CK(clk), .Q(
        fir_data[508]) );
  DFFTRX1 fir_data_reg_0__11_ ( .D(data[11]), .RN(n56), .CK(clk), .Q(
        fir_data[507]) );
  DFFTRX1 fir_data_reg_0__10_ ( .D(data[10]), .RN(n56), .CK(clk), .Q(
        fir_data[506]) );
  DFFTRX1 fir_data_reg_0__9_ ( .D(data[9]), .RN(n56), .CK(clk), .Q(
        fir_data[505]) );
  DFFTRX1 fir_data_reg_0__8_ ( .D(data[8]), .RN(n56), .CK(clk), .Q(
        fir_data[504]) );
  DFFTRX1 fir_data_reg_0__7_ ( .D(data[7]), .RN(n56), .CK(clk), .Q(
        fir_data[503]) );
  DFFTRX1 fir_data_reg_0__6_ ( .D(data[6]), .RN(n56), .CK(clk), .Q(
        fir_data[502]) );
  DFFTRX1 fir_data_reg_0__5_ ( .D(data[5]), .RN(n56), .CK(clk), .Q(
        fir_data[501]) );
  DFFQX1 fir_data_reg_31__11_ ( .D(fir_data[27]), .CK(clk), .Q(fir_data[11])
         );
  DFFQX1 fir_data_reg_31__10_ ( .D(fir_data[26]), .CK(clk), .Q(fir_data[10])
         );
  DFFQX1 fir_data_reg_31__9_ ( .D(fir_data[25]), .CK(clk), .Q(fir_data[9]) );
  DFFQX1 fir_data_reg_31__8_ ( .D(fir_data[24]), .CK(clk), .Q(fir_data[8]) );
  DFFQX1 fir_data_reg_31__7_ ( .D(fir_data[23]), .CK(clk), .Q(fir_data[7]) );
  DFFQX1 fir_data_reg_31__6_ ( .D(fir_data[22]), .CK(clk), .Q(fir_data[6]) );
  DFFQX1 fir_data_reg_31__5_ ( .D(fir_data[21]), .CK(clk), .Q(fir_data[5]) );
  DFFQX1 fir_data_reg_31__4_ ( .D(fir_data[20]), .CK(clk), .Q(fir_data[4]) );
  DFFQX1 temp_mul_add_fir_reg_1__31_ ( .D(mul_add_fir[456]), .CK(clk), .Q(
        temp_mul_add_fir[479]) );
  DFFQX1 temp_mul_add_fir_reg_1__30_ ( .D(mul_add_fir[455]), .CK(clk), .Q(
        temp_mul_add_fir[478]) );
  DFFQX1 temp_mul_add_fir_reg_1__29_ ( .D(mul_add_fir[454]), .CK(clk), .Q(
        temp_mul_add_fir[477]) );
  DFFQX1 temp_mul_add_fir_reg_1__28_ ( .D(mul_add_fir[453]), .CK(clk), .Q(
        temp_mul_add_fir[476]) );
  DFFQX1 temp_mul_add_fir_reg_3__31_ ( .D(mul_add_fir[393]), .CK(clk), .Q(
        temp_mul_add_fir[415]) );
  DFFQX1 temp_mul_add_fir_reg_3__30_ ( .D(mul_add_fir[392]), .CK(clk), .Q(
        temp_mul_add_fir[414]) );
  DFFQX1 temp_mul_add_fir_reg_3__29_ ( .D(mul_add_fir[391]), .CK(clk), .Q(
        temp_mul_add_fir[413]) );
  DFFQX1 temp_mul_add_fir_reg_3__28_ ( .D(mul_add_fir[390]), .CK(clk), .Q(
        temp_mul_add_fir[412]) );
  DFFQX1 temp_mul_add_fir_reg_5__31_ ( .D(mul_add_fir[329]), .CK(clk), .Q(
        temp_mul_add_fir[351]) );
  DFFQX1 temp_mul_add_fir_reg_5__30_ ( .D(mul_add_fir[328]), .CK(clk), .Q(
        temp_mul_add_fir[350]) );
  DFFQX1 temp_mul_add_fir_reg_5__29_ ( .D(mul_add_fir[327]), .CK(clk), .Q(
        temp_mul_add_fir[349]) );
  DFFQX1 temp_mul_add_fir_reg_5__28_ ( .D(mul_add_fir[326]), .CK(clk), .Q(
        temp_mul_add_fir[348]) );
  DFFQX1 temp_mul_add_fir_reg_7__31_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[287]) );
  DFFQX1 temp_mul_add_fir_reg_7__30_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[286]) );
  DFFQX1 temp_mul_add_fir_reg_7__29_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[285]) );
  DFFQX1 temp_mul_add_fir_reg_7__28_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[284]) );
  DFFQX1 temp_mul_add_fir_reg_9__31_ ( .D(mul_add_fir[215]), .CK(clk), .Q(
        temp_mul_add_fir[223]) );
  DFFQX1 temp_mul_add_fir_reg_9__30_ ( .D(mul_add_fir[214]), .CK(clk), .Q(
        temp_mul_add_fir[222]) );
  DFFQX1 temp_mul_add_fir_reg_9__29_ ( .D(mul_add_fir[213]), .CK(clk), .Q(
        temp_mul_add_fir[221]) );
  DFFQX1 temp_mul_add_fir_reg_9__28_ ( .D(mul_add_fir[212]), .CK(clk), .Q(
        temp_mul_add_fir[220]) );
  DFFQX1 temp_mul_add_fir_reg_11__31_ ( .D(mul_add_fir[153]), .CK(clk), .Q(
        temp_mul_add_fir[159]) );
  DFFQX1 temp_mul_add_fir_reg_11__30_ ( .D(mul_add_fir[152]), .CK(clk), .Q(
        temp_mul_add_fir[158]) );
  DFFQX1 temp_mul_add_fir_reg_11__29_ ( .D(mul_add_fir[151]), .CK(clk), .Q(
        temp_mul_add_fir[157]) );
  DFFQX1 temp_mul_add_fir_reg_11__28_ ( .D(mul_add_fir[150]), .CK(clk), .Q(
        temp_mul_add_fir[156]) );
  DFFQX1 temp_mul_add_fir_reg_13__31_ ( .D(mul_add_fir[92]), .CK(clk), .Q(
        temp_mul_add_fir[95]) );
  DFFQX1 temp_mul_add_fir_reg_13__30_ ( .D(mul_add_fir[91]), .CK(clk), .Q(
        temp_mul_add_fir[94]) );
  DFFQX1 temp_mul_add_fir_reg_13__29_ ( .D(mul_add_fir[90]), .CK(clk), .Q(
        temp_mul_add_fir[93]) );
  DFFQX1 temp_mul_add_fir_reg_13__28_ ( .D(mul_add_fir[89]), .CK(clk), .Q(
        temp_mul_add_fir[92]) );
  DFFQX1 temp_mul_add_fir_reg_15__31_ ( .D(mul_add_fir[31]), .CK(clk), .Q(
        temp_mul_add_fir[31]) );
  DFFQX1 temp_mul_add_fir_reg_15__30_ ( .D(mul_add_fir[30]), .CK(clk), .Q(
        temp_mul_add_fir[30]) );
  DFFQX1 temp_mul_add_fir_reg_15__29_ ( .D(mul_add_fir[29]), .CK(clk), .Q(
        temp_mul_add_fir[29]) );
  DFFQX1 temp_mul_add_fir_reg_15__28_ ( .D(mul_add_fir[28]), .CK(clk), .Q(
        temp_mul_add_fir[28]) );
  DFFQX1 temp_add_fir_reg_7__15_ ( .D(add_fir[143]), .CK(clk), .Q(
        temp_add_fir[140]) );
  DFFQX1 fir_data_reg_16__11_ ( .D(fir_data[267]), .CK(clk), .Q(fir_data[251])
         );
  DFFQX1 fir_data_reg_16__10_ ( .D(fir_data[266]), .CK(clk), .Q(fir_data[250])
         );
  DFFQX1 fir_data_reg_16__9_ ( .D(fir_data[265]), .CK(clk), .Q(fir_data[249])
         );
  DFFQX1 fir_data_reg_16__8_ ( .D(fir_data[264]), .CK(clk), .Q(fir_data[248])
         );
  DFFQX1 fir_data_reg_16__7_ ( .D(fir_data[263]), .CK(clk), .Q(fir_data[247])
         );
  DFFQX1 fir_data_reg_16__6_ ( .D(fir_data[262]), .CK(clk), .Q(fir_data[246])
         );
  DFFQX1 fir_data_reg_16__5_ ( .D(fir_data[261]), .CK(clk), .Q(fir_data[245])
         );
  DFFQX1 fir_data_reg_16__4_ ( .D(fir_data[260]), .CK(clk), .Q(fir_data[244])
         );
  DFFQX1 fir_data_reg_17__11_ ( .D(fir_data[251]), .CK(clk), .Q(fir_data[235])
         );
  DFFQX1 fir_data_reg_17__10_ ( .D(fir_data[250]), .CK(clk), .Q(fir_data[234])
         );
  DFFQX1 fir_data_reg_17__9_ ( .D(fir_data[249]), .CK(clk), .Q(fir_data[233])
         );
  DFFQX1 fir_data_reg_17__8_ ( .D(fir_data[248]), .CK(clk), .Q(fir_data[232])
         );
  DFFQX1 fir_data_reg_17__7_ ( .D(fir_data[247]), .CK(clk), .Q(fir_data[231])
         );
  DFFQX1 fir_data_reg_17__6_ ( .D(fir_data[246]), .CK(clk), .Q(fir_data[230])
         );
  DFFQX1 fir_data_reg_17__5_ ( .D(fir_data[245]), .CK(clk), .Q(fir_data[229])
         );
  DFFQX1 fir_data_reg_17__4_ ( .D(fir_data[244]), .CK(clk), .Q(fir_data[228])
         );
  DFFQX1 fir_data_reg_18__11_ ( .D(fir_data[235]), .CK(clk), .Q(fir_data[219])
         );
  DFFQX1 fir_data_reg_18__10_ ( .D(fir_data[234]), .CK(clk), .Q(fir_data[218])
         );
  DFFQX1 fir_data_reg_18__9_ ( .D(fir_data[233]), .CK(clk), .Q(fir_data[217])
         );
  DFFQX1 fir_data_reg_18__8_ ( .D(fir_data[232]), .CK(clk), .Q(fir_data[216])
         );
  DFFQX1 fir_data_reg_18__7_ ( .D(fir_data[231]), .CK(clk), .Q(fir_data[215])
         );
  DFFQX1 fir_data_reg_18__6_ ( .D(fir_data[230]), .CK(clk), .Q(fir_data[214])
         );
  DFFQX1 fir_data_reg_18__5_ ( .D(fir_data[229]), .CK(clk), .Q(fir_data[213])
         );
  DFFQX1 fir_data_reg_18__4_ ( .D(fir_data[228]), .CK(clk), .Q(fir_data[212])
         );
  DFFQX1 fir_data_reg_19__11_ ( .D(fir_data[219]), .CK(clk), .Q(fir_data[203])
         );
  DFFQX1 fir_data_reg_19__10_ ( .D(fir_data[218]), .CK(clk), .Q(fir_data[202])
         );
  DFFQX1 fir_data_reg_19__9_ ( .D(fir_data[217]), .CK(clk), .Q(fir_data[201])
         );
  DFFQX1 fir_data_reg_19__8_ ( .D(fir_data[216]), .CK(clk), .Q(fir_data[200])
         );
  DFFQX1 fir_data_reg_19__7_ ( .D(fir_data[215]), .CK(clk), .Q(fir_data[199])
         );
  DFFQX1 fir_data_reg_19__6_ ( .D(fir_data[214]), .CK(clk), .Q(fir_data[198])
         );
  DFFQX1 fir_data_reg_19__5_ ( .D(fir_data[213]), .CK(clk), .Q(fir_data[197])
         );
  DFFQX1 fir_data_reg_19__4_ ( .D(fir_data[212]), .CK(clk), .Q(fir_data[196])
         );
  DFFQX1 fir_data_reg_20__11_ ( .D(fir_data[203]), .CK(clk), .Q(fir_data[187])
         );
  DFFQX1 fir_data_reg_20__10_ ( .D(fir_data[202]), .CK(clk), .Q(fir_data[186])
         );
  DFFQX1 fir_data_reg_20__9_ ( .D(fir_data[201]), .CK(clk), .Q(fir_data[185])
         );
  DFFQX1 fir_data_reg_20__8_ ( .D(fir_data[200]), .CK(clk), .Q(fir_data[184])
         );
  DFFQX1 fir_data_reg_20__7_ ( .D(fir_data[199]), .CK(clk), .Q(fir_data[183])
         );
  DFFQX1 fir_data_reg_20__6_ ( .D(fir_data[198]), .CK(clk), .Q(fir_data[182])
         );
  DFFQX1 fir_data_reg_20__5_ ( .D(fir_data[197]), .CK(clk), .Q(fir_data[181])
         );
  DFFQX1 fir_data_reg_20__4_ ( .D(fir_data[196]), .CK(clk), .Q(fir_data[180])
         );
  DFFQX1 fir_data_reg_21__11_ ( .D(fir_data[187]), .CK(clk), .Q(fir_data[171])
         );
  DFFQX1 fir_data_reg_21__10_ ( .D(fir_data[186]), .CK(clk), .Q(fir_data[170])
         );
  DFFQX1 fir_data_reg_21__9_ ( .D(fir_data[185]), .CK(clk), .Q(fir_data[169])
         );
  DFFQX1 fir_data_reg_21__8_ ( .D(fir_data[184]), .CK(clk), .Q(fir_data[168])
         );
  DFFQX1 fir_data_reg_21__7_ ( .D(fir_data[183]), .CK(clk), .Q(fir_data[167])
         );
  DFFQX1 fir_data_reg_21__6_ ( .D(fir_data[182]), .CK(clk), .Q(fir_data[166])
         );
  DFFQX1 fir_data_reg_21__5_ ( .D(fir_data[181]), .CK(clk), .Q(fir_data[165])
         );
  DFFQX1 fir_data_reg_21__4_ ( .D(fir_data[180]), .CK(clk), .Q(fir_data[164])
         );
  DFFQX1 fir_data_reg_22__11_ ( .D(fir_data[171]), .CK(clk), .Q(fir_data[155])
         );
  DFFQX1 fir_data_reg_22__10_ ( .D(fir_data[170]), .CK(clk), .Q(fir_data[154])
         );
  DFFQX1 fir_data_reg_22__9_ ( .D(fir_data[169]), .CK(clk), .Q(fir_data[153])
         );
  DFFQX1 fir_data_reg_22__8_ ( .D(fir_data[168]), .CK(clk), .Q(fir_data[152])
         );
  DFFQX1 fir_data_reg_22__7_ ( .D(fir_data[167]), .CK(clk), .Q(fir_data[151])
         );
  DFFQX1 fir_data_reg_22__6_ ( .D(fir_data[166]), .CK(clk), .Q(fir_data[150])
         );
  DFFQX1 fir_data_reg_22__5_ ( .D(fir_data[165]), .CK(clk), .Q(fir_data[149])
         );
  DFFQX1 fir_data_reg_22__4_ ( .D(fir_data[164]), .CK(clk), .Q(fir_data[148])
         );
  DFFQX1 fir_data_reg_23__11_ ( .D(fir_data[155]), .CK(clk), .Q(fir_data[139])
         );
  DFFQX1 fir_data_reg_23__10_ ( .D(fir_data[154]), .CK(clk), .Q(fir_data[138])
         );
  DFFQX1 fir_data_reg_23__9_ ( .D(fir_data[153]), .CK(clk), .Q(fir_data[137])
         );
  DFFQX1 fir_data_reg_23__8_ ( .D(fir_data[152]), .CK(clk), .Q(fir_data[136])
         );
  DFFQX1 fir_data_reg_23__7_ ( .D(fir_data[151]), .CK(clk), .Q(fir_data[135])
         );
  DFFQX1 fir_data_reg_23__6_ ( .D(fir_data[150]), .CK(clk), .Q(fir_data[134])
         );
  DFFQX1 fir_data_reg_23__5_ ( .D(fir_data[149]), .CK(clk), .Q(fir_data[133])
         );
  DFFQX1 fir_data_reg_23__4_ ( .D(fir_data[148]), .CK(clk), .Q(fir_data[132])
         );
  DFFQX1 fir_data_reg_24__11_ ( .D(fir_data[139]), .CK(clk), .Q(fir_data[123])
         );
  DFFQX1 fir_data_reg_24__10_ ( .D(fir_data[138]), .CK(clk), .Q(fir_data[122])
         );
  DFFQX1 fir_data_reg_24__9_ ( .D(fir_data[137]), .CK(clk), .Q(fir_data[121])
         );
  DFFQX1 fir_data_reg_24__8_ ( .D(fir_data[136]), .CK(clk), .Q(fir_data[120])
         );
  DFFQX1 fir_data_reg_24__7_ ( .D(fir_data[135]), .CK(clk), .Q(fir_data[119])
         );
  DFFQX1 fir_data_reg_24__6_ ( .D(fir_data[134]), .CK(clk), .Q(fir_data[118])
         );
  DFFQX1 fir_data_reg_24__5_ ( .D(fir_data[133]), .CK(clk), .Q(fir_data[117])
         );
  DFFQX1 fir_data_reg_24__4_ ( .D(fir_data[132]), .CK(clk), .Q(fir_data[116])
         );
  DFFQX1 fir_data_reg_25__11_ ( .D(fir_data[123]), .CK(clk), .Q(fir_data[107])
         );
  DFFQX1 fir_data_reg_25__10_ ( .D(fir_data[122]), .CK(clk), .Q(fir_data[106])
         );
  DFFQX1 fir_data_reg_25__9_ ( .D(fir_data[121]), .CK(clk), .Q(fir_data[105])
         );
  DFFQX1 fir_data_reg_25__8_ ( .D(fir_data[120]), .CK(clk), .Q(fir_data[104])
         );
  DFFQX1 fir_data_reg_25__7_ ( .D(fir_data[119]), .CK(clk), .Q(fir_data[103])
         );
  DFFQX1 fir_data_reg_25__6_ ( .D(fir_data[118]), .CK(clk), .Q(fir_data[102])
         );
  DFFQX1 fir_data_reg_25__5_ ( .D(fir_data[117]), .CK(clk), .Q(fir_data[101])
         );
  DFFQX1 fir_data_reg_25__4_ ( .D(fir_data[116]), .CK(clk), .Q(fir_data[100])
         );
  DFFQX1 fir_data_reg_26__11_ ( .D(fir_data[107]), .CK(clk), .Q(fir_data[91])
         );
  DFFQX1 fir_data_reg_26__10_ ( .D(fir_data[106]), .CK(clk), .Q(fir_data[90])
         );
  DFFQX1 fir_data_reg_26__9_ ( .D(fir_data[105]), .CK(clk), .Q(fir_data[89])
         );
  DFFQX1 fir_data_reg_26__8_ ( .D(fir_data[104]), .CK(clk), .Q(fir_data[88])
         );
  DFFQX1 fir_data_reg_26__7_ ( .D(fir_data[103]), .CK(clk), .Q(fir_data[87])
         );
  DFFQX1 fir_data_reg_26__6_ ( .D(fir_data[102]), .CK(clk), .Q(fir_data[86])
         );
  DFFQX1 fir_data_reg_26__5_ ( .D(fir_data[101]), .CK(clk), .Q(fir_data[85])
         );
  DFFQX1 fir_data_reg_26__4_ ( .D(fir_data[100]), .CK(clk), .Q(fir_data[84])
         );
  DFFQX1 fir_data_reg_27__11_ ( .D(fir_data[91]), .CK(clk), .Q(fir_data[75])
         );
  DFFQX1 fir_data_reg_27__10_ ( .D(fir_data[90]), .CK(clk), .Q(fir_data[74])
         );
  DFFQX1 fir_data_reg_27__9_ ( .D(fir_data[89]), .CK(clk), .Q(fir_data[73]) );
  DFFQX1 fir_data_reg_27__8_ ( .D(fir_data[88]), .CK(clk), .Q(fir_data[72]) );
  DFFQX1 fir_data_reg_27__7_ ( .D(fir_data[87]), .CK(clk), .Q(fir_data[71]) );
  DFFQX1 fir_data_reg_27__6_ ( .D(fir_data[86]), .CK(clk), .Q(fir_data[70]) );
  DFFQX1 fir_data_reg_27__5_ ( .D(fir_data[85]), .CK(clk), .Q(fir_data[69]) );
  DFFQX1 fir_data_reg_27__4_ ( .D(fir_data[84]), .CK(clk), .Q(fir_data[68]) );
  DFFQX1 fir_data_reg_28__11_ ( .D(fir_data[75]), .CK(clk), .Q(fir_data[59])
         );
  DFFQX1 fir_data_reg_28__10_ ( .D(fir_data[74]), .CK(clk), .Q(fir_data[58])
         );
  DFFQX1 fir_data_reg_28__9_ ( .D(fir_data[73]), .CK(clk), .Q(fir_data[57]) );
  DFFQX1 fir_data_reg_28__8_ ( .D(fir_data[72]), .CK(clk), .Q(fir_data[56]) );
  DFFQX1 fir_data_reg_28__7_ ( .D(fir_data[71]), .CK(clk), .Q(fir_data[55]) );
  DFFQX1 fir_data_reg_28__6_ ( .D(fir_data[70]), .CK(clk), .Q(fir_data[54]) );
  DFFQX1 fir_data_reg_28__5_ ( .D(fir_data[69]), .CK(clk), .Q(fir_data[53]) );
  DFFQX1 fir_data_reg_28__4_ ( .D(fir_data[68]), .CK(clk), .Q(fir_data[52]) );
  DFFQX1 fir_data_reg_29__11_ ( .D(fir_data[59]), .CK(clk), .Q(fir_data[43])
         );
  DFFQX1 fir_data_reg_29__10_ ( .D(fir_data[58]), .CK(clk), .Q(fir_data[42])
         );
  DFFQX1 fir_data_reg_29__9_ ( .D(fir_data[57]), .CK(clk), .Q(fir_data[41]) );
  DFFQX1 fir_data_reg_29__8_ ( .D(fir_data[56]), .CK(clk), .Q(fir_data[40]) );
  DFFQX1 fir_data_reg_29__7_ ( .D(fir_data[55]), .CK(clk), .Q(fir_data[39]) );
  DFFQX1 fir_data_reg_29__6_ ( .D(fir_data[54]), .CK(clk), .Q(fir_data[38]) );
  DFFQX1 fir_data_reg_29__5_ ( .D(fir_data[53]), .CK(clk), .Q(fir_data[37]) );
  DFFQX1 fir_data_reg_29__4_ ( .D(fir_data[52]), .CK(clk), .Q(fir_data[36]) );
  DFFQX1 fir_data_reg_30__11_ ( .D(fir_data[43]), .CK(clk), .Q(fir_data[27])
         );
  DFFQX1 fir_data_reg_30__10_ ( .D(fir_data[42]), .CK(clk), .Q(fir_data[26])
         );
  DFFQX1 fir_data_reg_30__9_ ( .D(fir_data[41]), .CK(clk), .Q(fir_data[25]) );
  DFFQX1 fir_data_reg_30__8_ ( .D(fir_data[40]), .CK(clk), .Q(fir_data[24]) );
  DFFQX1 fir_data_reg_30__7_ ( .D(fir_data[39]), .CK(clk), .Q(fir_data[23]) );
  DFFQX1 fir_data_reg_30__6_ ( .D(fir_data[38]), .CK(clk), .Q(fir_data[22]) );
  DFFQX1 fir_data_reg_30__5_ ( .D(fir_data[37]), .CK(clk), .Q(fir_data[21]) );
  DFFQX1 fir_data_reg_30__4_ ( .D(fir_data[36]), .CK(clk), .Q(fir_data[20]) );
  DFFQX1 temp_mul_add_fir_reg_0__27_ ( .D(mul_add_fir[483]), .CK(clk), .Q(
        temp_mul_add_fir[507]) );
  DFFQX1 temp_mul_add_fir_reg_0__26_ ( .D(mul_add_fir[482]), .CK(clk), .Q(
        temp_mul_add_fir[506]) );
  DFFQX1 temp_mul_add_fir_reg_0__25_ ( .D(mul_add_fir[481]), .CK(clk), .Q(
        temp_mul_add_fir[505]) );
  DFFQX1 temp_mul_add_fir_reg_0__24_ ( .D(mul_add_fir[480]), .CK(clk), .Q(
        temp_mul_add_fir[504]) );
  DFFQX1 temp_mul_add_fir_reg_0__23_ ( .D(mul_add_fir[479]), .CK(clk), .Q(
        temp_mul_add_fir[503]) );
  DFFQX1 temp_mul_add_fir_reg_0__22_ ( .D(mul_add_fir[478]), .CK(clk), .Q(
        temp_mul_add_fir[502]) );
  DFFQX1 temp_mul_add_fir_reg_0__21_ ( .D(mul_add_fir[477]), .CK(clk), .Q(
        temp_mul_add_fir[501]) );
  DFFQX1 temp_mul_add_fir_reg_2__27_ ( .D(mul_add_fir[421]), .CK(clk), .Q(
        temp_mul_add_fir[443]) );
  DFFQX1 temp_mul_add_fir_reg_2__26_ ( .D(mul_add_fir[420]), .CK(clk), .Q(
        temp_mul_add_fir[442]) );
  DFFQX1 temp_mul_add_fir_reg_2__25_ ( .D(mul_add_fir[419]), .CK(clk), .Q(
        temp_mul_add_fir[441]) );
  DFFQX1 temp_mul_add_fir_reg_2__24_ ( .D(mul_add_fir[418]), .CK(clk), .Q(
        temp_mul_add_fir[440]) );
  DFFQX1 temp_mul_add_fir_reg_2__23_ ( .D(mul_add_fir[417]), .CK(clk), .Q(
        temp_mul_add_fir[439]) );
  DFFQX1 temp_mul_add_fir_reg_2__22_ ( .D(mul_add_fir[416]), .CK(clk), .Q(
        temp_mul_add_fir[438]) );
  DFFQX1 temp_mul_add_fir_reg_2__21_ ( .D(mul_add_fir[415]), .CK(clk), .Q(
        temp_mul_add_fir[437]) );
  DFFQX1 temp_mul_add_fir_reg_2__20_ ( .D(mul_add_fir[414]), .CK(clk), .Q(
        temp_mul_add_fir[436]) );
  DFFQX1 temp_mul_add_fir_reg_4__27_ ( .D(mul_add_fir[357]), .CK(clk), .Q(
        temp_mul_add_fir[379]) );
  DFFQX1 temp_mul_add_fir_reg_4__26_ ( .D(mul_add_fir[356]), .CK(clk), .Q(
        temp_mul_add_fir[378]) );
  DFFQX1 temp_mul_add_fir_reg_4__25_ ( .D(mul_add_fir[355]), .CK(clk), .Q(
        temp_mul_add_fir[377]) );
  DFFQX1 temp_mul_add_fir_reg_4__24_ ( .D(mul_add_fir[354]), .CK(clk), .Q(
        temp_mul_add_fir[376]) );
  DFFQX1 temp_mul_add_fir_reg_4__23_ ( .D(mul_add_fir[353]), .CK(clk), .Q(
        temp_mul_add_fir[375]) );
  DFFQX1 temp_mul_add_fir_reg_4__22_ ( .D(mul_add_fir[352]), .CK(clk), .Q(
        temp_mul_add_fir[374]) );
  DFFQX1 temp_mul_add_fir_reg_4__21_ ( .D(mul_add_fir[351]), .CK(clk), .Q(
        temp_mul_add_fir[373]) );
  DFFQX1 temp_mul_add_fir_reg_4__20_ ( .D(mul_add_fir[350]), .CK(clk), .Q(
        temp_mul_add_fir[372]) );
  DFFQX1 temp_mul_add_fir_reg_6__27_ ( .D(mul_add_fir[294]), .CK(clk), .Q(
        temp_mul_add_fir[315]) );
  DFFQX1 temp_mul_add_fir_reg_6__26_ ( .D(mul_add_fir[293]), .CK(clk), .Q(
        temp_mul_add_fir[314]) );
  DFFQX1 temp_mul_add_fir_reg_6__25_ ( .D(mul_add_fir[292]), .CK(clk), .Q(
        temp_mul_add_fir[313]) );
  DFFQX1 temp_mul_add_fir_reg_6__24_ ( .D(mul_add_fir[291]), .CK(clk), .Q(
        temp_mul_add_fir[312]) );
  DFFQX1 temp_mul_add_fir_reg_6__23_ ( .D(mul_add_fir[290]), .CK(clk), .Q(
        temp_mul_add_fir[311]) );
  DFFQX1 temp_mul_add_fir_reg_6__22_ ( .D(mul_add_fir[289]), .CK(clk), .Q(
        temp_mul_add_fir[310]) );
  DFFQX1 temp_mul_add_fir_reg_6__21_ ( .D(mul_add_fir[288]), .CK(clk), .Q(
        temp_mul_add_fir[309]) );
  DFFQX1 temp_mul_add_fir_reg_6__20_ ( .D(mul_add_fir[287]), .CK(clk), .Q(
        temp_mul_add_fir[308]) );
  DFFQX1 temp_mul_add_fir_reg_8__27_ ( .D(mul_add_fir[243]), .CK(clk), .Q(
        temp_mul_add_fir[251]) );
  DFFQX1 temp_mul_add_fir_reg_8__26_ ( .D(mul_add_fir[242]), .CK(clk), .Q(
        temp_mul_add_fir[250]) );
  DFFQX1 temp_mul_add_fir_reg_8__25_ ( .D(mul_add_fir[241]), .CK(clk), .Q(
        temp_mul_add_fir[249]) );
  DFFQX1 temp_mul_add_fir_reg_8__24_ ( .D(mul_add_fir[240]), .CK(clk), .Q(
        temp_mul_add_fir[248]) );
  DFFQX1 temp_mul_add_fir_reg_8__23_ ( .D(mul_add_fir[239]), .CK(clk), .Q(
        temp_mul_add_fir[247]) );
  DFFQX1 temp_mul_add_fir_reg_8__22_ ( .D(mul_add_fir[238]), .CK(clk), .Q(
        temp_mul_add_fir[246]) );
  DFFQX1 temp_mul_add_fir_reg_8__21_ ( .D(mul_add_fir[237]), .CK(clk), .Q(
        temp_mul_add_fir[245]) );
  DFFQX1 temp_mul_add_fir_reg_8__20_ ( .D(mul_add_fir[236]), .CK(clk), .Q(
        temp_mul_add_fir[244]) );
  DFFQX1 temp_mul_add_fir_reg_10__27_ ( .D(mul_add_fir[180]), .CK(clk), .Q(
        temp_mul_add_fir[187]) );
  DFFQX1 temp_mul_add_fir_reg_10__26_ ( .D(mul_add_fir[179]), .CK(clk), .Q(
        temp_mul_add_fir[186]) );
  DFFQX1 temp_mul_add_fir_reg_10__25_ ( .D(mul_add_fir[178]), .CK(clk), .Q(
        temp_mul_add_fir[185]) );
  DFFQX1 temp_mul_add_fir_reg_10__24_ ( .D(mul_add_fir[177]), .CK(clk), .Q(
        temp_mul_add_fir[184]) );
  DFFQX1 temp_mul_add_fir_reg_10__23_ ( .D(mul_add_fir[176]), .CK(clk), .Q(
        temp_mul_add_fir[183]) );
  DFFQX1 temp_mul_add_fir_reg_10__22_ ( .D(mul_add_fir[175]), .CK(clk), .Q(
        temp_mul_add_fir[182]) );
  DFFQX1 temp_mul_add_fir_reg_10__21_ ( .D(mul_add_fir[174]), .CK(clk), .Q(
        temp_mul_add_fir[181]) );
  DFFQX1 temp_mul_add_fir_reg_10__20_ ( .D(mul_add_fir[173]), .CK(clk), .Q(
        temp_mul_add_fir[180]) );
  DFFQX1 temp_mul_add_fir_reg_12__27_ ( .D(mul_add_fir[119]), .CK(clk), .Q(
        temp_mul_add_fir[123]) );
  DFFQX1 temp_mul_add_fir_reg_12__26_ ( .D(mul_add_fir[118]), .CK(clk), .Q(
        temp_mul_add_fir[122]) );
  DFFQX1 temp_mul_add_fir_reg_12__25_ ( .D(mul_add_fir[117]), .CK(clk), .Q(
        temp_mul_add_fir[121]) );
  DFFQX1 temp_mul_add_fir_reg_12__24_ ( .D(mul_add_fir[116]), .CK(clk), .Q(
        temp_mul_add_fir[120]) );
  DFFQX1 temp_mul_add_fir_reg_12__23_ ( .D(mul_add_fir[115]), .CK(clk), .Q(
        temp_mul_add_fir[119]) );
  DFFQX1 temp_mul_add_fir_reg_12__22_ ( .D(mul_add_fir[114]), .CK(clk), .Q(
        temp_mul_add_fir[118]) );
  DFFQX1 temp_mul_add_fir_reg_12__21_ ( .D(mul_add_fir[113]), .CK(clk), .Q(
        temp_mul_add_fir[117]) );
  DFFQX1 temp_mul_add_fir_reg_12__20_ ( .D(mul_add_fir[112]), .CK(clk), .Q(
        temp_mul_add_fir[116]) );
  DFFQX1 temp_mul_add_fir_reg_14__27_ ( .D(mul_add_fir[58]), .CK(clk), .Q(
        temp_mul_add_fir[59]) );
  DFFQX1 temp_mul_add_fir_reg_14__26_ ( .D(mul_add_fir[57]), .CK(clk), .Q(
        temp_mul_add_fir[58]) );
  DFFQX1 temp_mul_add_fir_reg_14__25_ ( .D(mul_add_fir[56]), .CK(clk), .Q(
        temp_mul_add_fir[57]) );
  DFFQX1 temp_mul_add_fir_reg_14__24_ ( .D(mul_add_fir[55]), .CK(clk), .Q(
        temp_mul_add_fir[56]) );
  DFFQX1 temp_mul_add_fir_reg_14__23_ ( .D(mul_add_fir[54]), .CK(clk), .Q(
        temp_mul_add_fir[55]) );
  DFFQX1 temp_mul_add_fir_reg_14__22_ ( .D(mul_add_fir[53]), .CK(clk), .Q(
        temp_mul_add_fir[54]) );
  DFFQX1 temp_mul_add_fir_reg_14__21_ ( .D(mul_add_fir[52]), .CK(clk), .Q(
        temp_mul_add_fir[53]) );
  DFFQX1 temp_mul_add_fir_reg_14__20_ ( .D(mul_add_fir[51]), .CK(clk), .Q(
        temp_mul_add_fir[52]) );
  DFFQX1 temp_add_fir_reg_7__12_ ( .D(add_fir[140]), .CK(clk), .Q(
        temp_add_fir[137]) );
  DFFQX1 fir_data_reg_1__3_ ( .D(fir_data[499]), .CK(clk), .Q(fir_data[483])
         );
  DFFQX1 fir_data_reg_1__2_ ( .D(fir_data[498]), .CK(clk), .Q(fir_data[482])
         );
  DFFQX1 fir_data_reg_1__1_ ( .D(fir_data[497]), .CK(clk), .Q(fir_data[481])
         );
  DFFQX1 fir_data_reg_2__3_ ( .D(fir_data[483]), .CK(clk), .Q(fir_data[467])
         );
  DFFQX1 fir_data_reg_2__2_ ( .D(fir_data[482]), .CK(clk), .Q(fir_data[466])
         );
  DFFQX1 fir_data_reg_2__1_ ( .D(fir_data[481]), .CK(clk), .Q(fir_data[465])
         );
  DFFQX1 fir_data_reg_3__3_ ( .D(fir_data[467]), .CK(clk), .Q(fir_data[451])
         );
  DFFQX1 fir_data_reg_3__2_ ( .D(fir_data[466]), .CK(clk), .Q(fir_data[450])
         );
  DFFQX1 fir_data_reg_3__1_ ( .D(fir_data[465]), .CK(clk), .Q(fir_data[449])
         );
  DFFQX1 fir_data_reg_4__3_ ( .D(fir_data[451]), .CK(clk), .Q(fir_data[435])
         );
  DFFQX1 fir_data_reg_4__2_ ( .D(fir_data[450]), .CK(clk), .Q(fir_data[434])
         );
  DFFQX1 fir_data_reg_4__1_ ( .D(fir_data[449]), .CK(clk), .Q(fir_data[433])
         );
  DFFQX1 fir_data_reg_5__3_ ( .D(fir_data[435]), .CK(clk), .Q(fir_data[419])
         );
  DFFQX1 fir_data_reg_5__2_ ( .D(fir_data[434]), .CK(clk), .Q(fir_data[418])
         );
  DFFQX1 fir_data_reg_5__1_ ( .D(fir_data[433]), .CK(clk), .Q(fir_data[417])
         );
  DFFQX1 fir_data_reg_6__3_ ( .D(fir_data[419]), .CK(clk), .Q(fir_data[403])
         );
  DFFQX1 fir_data_reg_6__2_ ( .D(fir_data[418]), .CK(clk), .Q(fir_data[402])
         );
  DFFQX1 fir_data_reg_6__1_ ( .D(fir_data[417]), .CK(clk), .Q(fir_data[401])
         );
  DFFQX1 fir_data_reg_7__3_ ( .D(fir_data[403]), .CK(clk), .Q(fir_data[387])
         );
  DFFQX1 fir_data_reg_7__2_ ( .D(fir_data[402]), .CK(clk), .Q(fir_data[386])
         );
  DFFQX1 fir_data_reg_7__1_ ( .D(fir_data[401]), .CK(clk), .Q(fir_data[385])
         );
  DFFQX1 fir_data_reg_8__3_ ( .D(fir_data[387]), .CK(clk), .Q(fir_data[371])
         );
  DFFQX1 fir_data_reg_8__2_ ( .D(fir_data[386]), .CK(clk), .Q(fir_data[370])
         );
  DFFQX1 fir_data_reg_8__1_ ( .D(fir_data[385]), .CK(clk), .Q(fir_data[369])
         );
  DFFQX1 fir_data_reg_9__3_ ( .D(fir_data[371]), .CK(clk), .Q(fir_data[355])
         );
  DFFQX1 fir_data_reg_9__2_ ( .D(fir_data[370]), .CK(clk), .Q(fir_data[354])
         );
  DFFQX1 fir_data_reg_9__1_ ( .D(fir_data[369]), .CK(clk), .Q(fir_data[353])
         );
  DFFQX1 fir_data_reg_10__3_ ( .D(fir_data[355]), .CK(clk), .Q(fir_data[339])
         );
  DFFQX1 fir_data_reg_10__2_ ( .D(fir_data[354]), .CK(clk), .Q(fir_data[338])
         );
  DFFQX1 fir_data_reg_10__1_ ( .D(fir_data[353]), .CK(clk), .Q(fir_data[337])
         );
  DFFQX1 fir_data_reg_11__3_ ( .D(fir_data[339]), .CK(clk), .Q(fir_data[323])
         );
  DFFQX1 fir_data_reg_11__2_ ( .D(fir_data[338]), .CK(clk), .Q(fir_data[322])
         );
  DFFQX1 fir_data_reg_11__1_ ( .D(fir_data[337]), .CK(clk), .Q(fir_data[321])
         );
  DFFQX1 fir_data_reg_12__3_ ( .D(fir_data[323]), .CK(clk), .Q(fir_data[307])
         );
  DFFQX1 fir_data_reg_12__2_ ( .D(fir_data[322]), .CK(clk), .Q(fir_data[306])
         );
  DFFQX1 fir_data_reg_12__1_ ( .D(fir_data[321]), .CK(clk), .Q(fir_data[305])
         );
  DFFQX1 fir_data_reg_13__3_ ( .D(fir_data[307]), .CK(clk), .Q(fir_data[291])
         );
  DFFQX1 fir_data_reg_13__2_ ( .D(fir_data[306]), .CK(clk), .Q(fir_data[290])
         );
  DFFQX1 fir_data_reg_13__1_ ( .D(fir_data[305]), .CK(clk), .Q(fir_data[289])
         );
  DFFQX1 fir_data_reg_14__3_ ( .D(fir_data[291]), .CK(clk), .Q(fir_data[275])
         );
  DFFQX1 fir_data_reg_14__2_ ( .D(fir_data[290]), .CK(clk), .Q(fir_data[274])
         );
  DFFQX1 fir_data_reg_14__1_ ( .D(fir_data[289]), .CK(clk), .Q(fir_data[273])
         );
  DFFQX1 fir_data_reg_15__3_ ( .D(fir_data[275]), .CK(clk), .Q(fir_data[259])
         );
  DFFQX1 fir_data_reg_15__2_ ( .D(fir_data[274]), .CK(clk), .Q(fir_data[258])
         );
  DFFQX1 fir_data_reg_15__1_ ( .D(fir_data[273]), .CK(clk), .Q(fir_data[257])
         );
  DFFTRX1 fir_data_reg_0__4_ ( .D(data[4]), .RN(n56), .CK(clk), .Q(
        fir_data[500]) );
  DFFTRX1 fir_data_reg_0__3_ ( .D(data[3]), .RN(n56), .CK(clk), .Q(
        fir_data[499]) );
  DFFTRX1 fir_data_reg_0__2_ ( .D(data[2]), .RN(n56), .CK(clk), .Q(
        fir_data[498]) );
  DFFTRX1 fir_data_reg_0__1_ ( .D(data[1]), .RN(n56), .CK(clk), .Q(
        fir_data[497]) );
  DFFQX1 fir_data_reg_31__0_ ( .D(fir_data[16]), .CK(clk), .Q(fir_data[0]) );
  DFFQX1 fir_data_reg_31__3_ ( .D(fir_data[19]), .CK(clk), .Q(fir_data[3]) );
  DFFQX1 fir_data_reg_31__2_ ( .D(fir_data[18]), .CK(clk), .Q(fir_data[2]) );
  DFFQX1 fir_data_reg_31__1_ ( .D(fir_data[17]), .CK(clk), .Q(fir_data[1]) );
  DFFQX1 temp_mul_add_fir_reg_1__27_ ( .D(mul_add_fir[452]), .CK(clk), .Q(
        temp_mul_add_fir[475]) );
  DFFQX1 temp_mul_add_fir_reg_1__26_ ( .D(mul_add_fir[451]), .CK(clk), .Q(
        temp_mul_add_fir[474]) );
  DFFQX1 temp_mul_add_fir_reg_1__25_ ( .D(mul_add_fir[450]), .CK(clk), .Q(
        temp_mul_add_fir[473]) );
  DFFQX1 temp_mul_add_fir_reg_1__24_ ( .D(mul_add_fir[449]), .CK(clk), .Q(
        temp_mul_add_fir[472]) );
  DFFQX1 temp_mul_add_fir_reg_1__23_ ( .D(mul_add_fir[448]), .CK(clk), .Q(
        temp_mul_add_fir[471]) );
  DFFQX1 temp_mul_add_fir_reg_1__22_ ( .D(mul_add_fir[447]), .CK(clk), .Q(
        temp_mul_add_fir[470]) );
  DFFQX1 temp_mul_add_fir_reg_1__21_ ( .D(mul_add_fir[446]), .CK(clk), .Q(
        temp_mul_add_fir[469]) );
  DFFQX1 temp_mul_add_fir_reg_1__20_ ( .D(mul_add_fir[445]), .CK(clk), .Q(
        temp_mul_add_fir[468]) );
  DFFQX1 temp_mul_add_fir_reg_3__27_ ( .D(mul_add_fir[389]), .CK(clk), .Q(
        temp_mul_add_fir[411]) );
  DFFQX1 temp_mul_add_fir_reg_3__26_ ( .D(mul_add_fir[388]), .CK(clk), .Q(
        temp_mul_add_fir[410]) );
  DFFQX1 temp_mul_add_fir_reg_3__25_ ( .D(mul_add_fir[387]), .CK(clk), .Q(
        temp_mul_add_fir[409]) );
  DFFQX1 temp_mul_add_fir_reg_3__24_ ( .D(mul_add_fir[386]), .CK(clk), .Q(
        temp_mul_add_fir[408]) );
  DFFQX1 temp_mul_add_fir_reg_3__23_ ( .D(mul_add_fir[385]), .CK(clk), .Q(
        temp_mul_add_fir[407]) );
  DFFQX1 temp_mul_add_fir_reg_3__22_ ( .D(mul_add_fir[384]), .CK(clk), .Q(
        temp_mul_add_fir[406]) );
  DFFQX1 temp_mul_add_fir_reg_3__21_ ( .D(mul_add_fir[383]), .CK(clk), .Q(
        temp_mul_add_fir[405]) );
  DFFQX1 temp_mul_add_fir_reg_3__20_ ( .D(mul_add_fir[382]), .CK(clk), .Q(
        temp_mul_add_fir[404]) );
  DFFQX1 temp_mul_add_fir_reg_5__27_ ( .D(mul_add_fir[325]), .CK(clk), .Q(
        temp_mul_add_fir[347]) );
  DFFQX1 temp_mul_add_fir_reg_5__26_ ( .D(mul_add_fir[324]), .CK(clk), .Q(
        temp_mul_add_fir[346]) );
  DFFQX1 temp_mul_add_fir_reg_5__25_ ( .D(mul_add_fir[323]), .CK(clk), .Q(
        temp_mul_add_fir[345]) );
  DFFQX1 temp_mul_add_fir_reg_5__24_ ( .D(mul_add_fir[322]), .CK(clk), .Q(
        temp_mul_add_fir[344]) );
  DFFQX1 temp_mul_add_fir_reg_5__23_ ( .D(mul_add_fir[321]), .CK(clk), .Q(
        temp_mul_add_fir[343]) );
  DFFQX1 temp_mul_add_fir_reg_5__22_ ( .D(mul_add_fir[320]), .CK(clk), .Q(
        temp_mul_add_fir[342]) );
  DFFQX1 temp_mul_add_fir_reg_5__21_ ( .D(mul_add_fir[319]), .CK(clk), .Q(
        temp_mul_add_fir[341]) );
  DFFQX1 temp_mul_add_fir_reg_5__20_ ( .D(mul_add_fir[318]), .CK(clk), .Q(
        temp_mul_add_fir[340]) );
  DFFQX1 temp_mul_add_fir_reg_7__27_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[283]) );
  DFFQX1 temp_mul_add_fir_reg_7__26_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[282]) );
  DFFQX1 temp_mul_add_fir_reg_7__25_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[281]) );
  DFFQX1 temp_mul_add_fir_reg_7__24_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[280]) );
  DFFQX1 temp_mul_add_fir_reg_7__23_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[279]) );
  DFFQX1 temp_mul_add_fir_reg_7__22_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[278]) );
  DFFQX1 temp_mul_add_fir_reg_7__21_ ( .D(n55), .CK(clk), .Q(
        temp_mul_add_fir[277]) );
  DFFQX1 temp_mul_add_fir_reg_7__20_ ( .D(mul_add_fir[266]), .CK(clk), .Q(
        temp_mul_add_fir[276]) );
  DFFQX1 temp_mul_add_fir_reg_9__27_ ( .D(mul_add_fir[211]), .CK(clk), .Q(
        temp_mul_add_fir[219]) );
  DFFQX1 temp_mul_add_fir_reg_9__26_ ( .D(mul_add_fir[210]), .CK(clk), .Q(
        temp_mul_add_fir[218]) );
  DFFQX1 temp_mul_add_fir_reg_9__25_ ( .D(mul_add_fir[209]), .CK(clk), .Q(
        temp_mul_add_fir[217]) );
  DFFQX1 temp_mul_add_fir_reg_9__24_ ( .D(mul_add_fir[208]), .CK(clk), .Q(
        temp_mul_add_fir[216]) );
  DFFQX1 temp_mul_add_fir_reg_9__23_ ( .D(mul_add_fir[207]), .CK(clk), .Q(
        temp_mul_add_fir[215]) );
  DFFQX1 temp_mul_add_fir_reg_9__22_ ( .D(mul_add_fir[206]), .CK(clk), .Q(
        temp_mul_add_fir[214]) );
  DFFQX1 temp_mul_add_fir_reg_9__21_ ( .D(mul_add_fir[205]), .CK(clk), .Q(
        temp_mul_add_fir[213]) );
  DFFQX1 temp_mul_add_fir_reg_9__20_ ( .D(mul_add_fir[204]), .CK(clk), .Q(
        temp_mul_add_fir[212]) );
  DFFQX1 temp_mul_add_fir_reg_11__27_ ( .D(mul_add_fir[149]), .CK(clk), .Q(
        temp_mul_add_fir[155]) );
  DFFQX1 temp_mul_add_fir_reg_11__26_ ( .D(mul_add_fir[148]), .CK(clk), .Q(
        temp_mul_add_fir[154]) );
  DFFQX1 temp_mul_add_fir_reg_11__25_ ( .D(mul_add_fir[147]), .CK(clk), .Q(
        temp_mul_add_fir[153]) );
  DFFQX1 temp_mul_add_fir_reg_11__24_ ( .D(mul_add_fir[146]), .CK(clk), .Q(
        temp_mul_add_fir[152]) );
  DFFQX1 temp_mul_add_fir_reg_11__23_ ( .D(mul_add_fir[145]), .CK(clk), .Q(
        temp_mul_add_fir[151]) );
  DFFQX1 temp_mul_add_fir_reg_11__22_ ( .D(mul_add_fir[144]), .CK(clk), .Q(
        temp_mul_add_fir[150]) );
  DFFQX1 temp_mul_add_fir_reg_11__21_ ( .D(mul_add_fir[143]), .CK(clk), .Q(
        temp_mul_add_fir[149]) );
  DFFQX1 temp_mul_add_fir_reg_11__20_ ( .D(mul_add_fir[142]), .CK(clk), .Q(
        temp_mul_add_fir[148]) );
  DFFQX1 temp_mul_add_fir_reg_13__27_ ( .D(mul_add_fir[88]), .CK(clk), .Q(
        temp_mul_add_fir[91]) );
  DFFQX1 temp_mul_add_fir_reg_13__26_ ( .D(mul_add_fir[87]), .CK(clk), .Q(
        temp_mul_add_fir[90]) );
  DFFQX1 temp_mul_add_fir_reg_13__25_ ( .D(mul_add_fir[86]), .CK(clk), .Q(
        temp_mul_add_fir[89]) );
  DFFQX1 temp_mul_add_fir_reg_13__24_ ( .D(mul_add_fir[85]), .CK(clk), .Q(
        temp_mul_add_fir[88]) );
  DFFQX1 temp_mul_add_fir_reg_13__23_ ( .D(mul_add_fir[84]), .CK(clk), .Q(
        temp_mul_add_fir[87]) );
  DFFQX1 temp_mul_add_fir_reg_13__22_ ( .D(mul_add_fir[83]), .CK(clk), .Q(
        temp_mul_add_fir[86]) );
  DFFQX1 temp_mul_add_fir_reg_13__21_ ( .D(mul_add_fir[82]), .CK(clk), .Q(
        temp_mul_add_fir[85]) );
  DFFQX1 temp_mul_add_fir_reg_13__20_ ( .D(mul_add_fir[81]), .CK(clk), .Q(
        temp_mul_add_fir[84]) );
  DFFQX1 temp_mul_add_fir_reg_15__27_ ( .D(mul_add_fir[27]), .CK(clk), .Q(
        temp_mul_add_fir[27]) );
  DFFQX1 temp_mul_add_fir_reg_15__26_ ( .D(mul_add_fir[26]), .CK(clk), .Q(
        temp_mul_add_fir[26]) );
  DFFQX1 temp_mul_add_fir_reg_15__25_ ( .D(mul_add_fir[25]), .CK(clk), .Q(
        temp_mul_add_fir[25]) );
  DFFQX1 temp_mul_add_fir_reg_15__24_ ( .D(mul_add_fir[24]), .CK(clk), .Q(
        temp_mul_add_fir[24]) );
  DFFQX1 temp_mul_add_fir_reg_15__23_ ( .D(mul_add_fir[23]), .CK(clk), .Q(
        temp_mul_add_fir[23]) );
  DFFQX1 temp_mul_add_fir_reg_15__22_ ( .D(mul_add_fir[22]), .CK(clk), .Q(
        temp_mul_add_fir[22]) );
  DFFQX1 temp_mul_add_fir_reg_15__21_ ( .D(mul_add_fir[21]), .CK(clk), .Q(
        temp_mul_add_fir[21]) );
  DFFQX1 temp_mul_add_fir_reg_15__20_ ( .D(mul_add_fir[20]), .CK(clk), .Q(
        temp_mul_add_fir[20]) );
  DFFQX1 temp_add_fir_reg_7__14_ ( .D(add_fir[142]), .CK(clk), .Q(
        temp_add_fir[139]) );
  DFFQX1 temp_add_fir_reg_7__13_ ( .D(add_fir[141]), .CK(clk), .Q(
        temp_add_fir[138]) );
  DFFQX1 fir_data_reg_16__0_ ( .D(fir_data[256]), .CK(clk), .Q(fir_data[240])
         );
  DFFQX1 fir_data_reg_17__0_ ( .D(fir_data[240]), .CK(clk), .Q(fir_data[224])
         );
  DFFQX1 fir_data_reg_18__0_ ( .D(fir_data[224]), .CK(clk), .Q(fir_data[208])
         );
  DFFQX1 fir_data_reg_19__0_ ( .D(fir_data[208]), .CK(clk), .Q(fir_data[192])
         );
  DFFQX1 fir_data_reg_20__0_ ( .D(fir_data[192]), .CK(clk), .Q(fir_data[176])
         );
  DFFQX1 fir_data_reg_21__0_ ( .D(fir_data[176]), .CK(clk), .Q(fir_data[160])
         );
  DFFQX1 fir_data_reg_22__0_ ( .D(fir_data[160]), .CK(clk), .Q(fir_data[144])
         );
  DFFQX1 fir_data_reg_23__0_ ( .D(fir_data[144]), .CK(clk), .Q(fir_data[128])
         );
  DFFQX1 fir_data_reg_24__0_ ( .D(fir_data[128]), .CK(clk), .Q(fir_data[112])
         );
  DFFQX1 fir_data_reg_25__0_ ( .D(fir_data[112]), .CK(clk), .Q(fir_data[96])
         );
  DFFQX1 fir_data_reg_26__0_ ( .D(fir_data[96]), .CK(clk), .Q(fir_data[80]) );
  DFFQX1 fir_data_reg_27__0_ ( .D(fir_data[80]), .CK(clk), .Q(fir_data[64]) );
  DFFQX1 fir_data_reg_28__0_ ( .D(fir_data[64]), .CK(clk), .Q(fir_data[48]) );
  DFFQX1 fir_data_reg_29__0_ ( .D(fir_data[48]), .CK(clk), .Q(fir_data[32]) );
  DFFQX1 fir_data_reg_30__0_ ( .D(fir_data[32]), .CK(clk), .Q(fir_data[16]) );
  DFFQX1 fir_data_reg_16__3_ ( .D(fir_data[259]), .CK(clk), .Q(fir_data[243])
         );
  DFFQX1 fir_data_reg_16__2_ ( .D(fir_data[258]), .CK(clk), .Q(fir_data[242])
         );
  DFFQX1 fir_data_reg_16__1_ ( .D(fir_data[257]), .CK(clk), .Q(fir_data[241])
         );
  DFFQX1 fir_data_reg_17__3_ ( .D(fir_data[243]), .CK(clk), .Q(fir_data[227])
         );
  DFFQX1 fir_data_reg_17__2_ ( .D(fir_data[242]), .CK(clk), .Q(fir_data[226])
         );
  DFFQX1 fir_data_reg_17__1_ ( .D(fir_data[241]), .CK(clk), .Q(fir_data[225])
         );
  DFFQX1 fir_data_reg_18__3_ ( .D(fir_data[227]), .CK(clk), .Q(fir_data[211])
         );
  DFFQX1 fir_data_reg_18__2_ ( .D(fir_data[226]), .CK(clk), .Q(fir_data[210])
         );
  DFFQX1 fir_data_reg_18__1_ ( .D(fir_data[225]), .CK(clk), .Q(fir_data[209])
         );
  DFFQX1 fir_data_reg_19__3_ ( .D(fir_data[211]), .CK(clk), .Q(fir_data[195])
         );
  DFFQX1 fir_data_reg_19__2_ ( .D(fir_data[210]), .CK(clk), .Q(fir_data[194])
         );
  DFFQX1 fir_data_reg_19__1_ ( .D(fir_data[209]), .CK(clk), .Q(fir_data[193])
         );
  DFFQX1 fir_data_reg_20__3_ ( .D(fir_data[195]), .CK(clk), .Q(fir_data[179])
         );
  DFFQX1 fir_data_reg_20__2_ ( .D(fir_data[194]), .CK(clk), .Q(fir_data[178])
         );
  DFFQX1 fir_data_reg_20__1_ ( .D(fir_data[193]), .CK(clk), .Q(fir_data[177])
         );
  DFFQX1 fir_data_reg_21__3_ ( .D(fir_data[179]), .CK(clk), .Q(fir_data[163])
         );
  DFFQX1 fir_data_reg_21__2_ ( .D(fir_data[178]), .CK(clk), .Q(fir_data[162])
         );
  DFFQX1 fir_data_reg_21__1_ ( .D(fir_data[177]), .CK(clk), .Q(fir_data[161])
         );
  DFFQX1 fir_data_reg_22__3_ ( .D(fir_data[163]), .CK(clk), .Q(fir_data[147])
         );
  DFFQX1 fir_data_reg_22__2_ ( .D(fir_data[162]), .CK(clk), .Q(fir_data[146])
         );
  DFFQX1 fir_data_reg_22__1_ ( .D(fir_data[161]), .CK(clk), .Q(fir_data[145])
         );
  DFFQX1 fir_data_reg_23__3_ ( .D(fir_data[147]), .CK(clk), .Q(fir_data[131])
         );
  DFFQX1 fir_data_reg_23__2_ ( .D(fir_data[146]), .CK(clk), .Q(fir_data[130])
         );
  DFFQX1 fir_data_reg_23__1_ ( .D(fir_data[145]), .CK(clk), .Q(fir_data[129])
         );
  DFFQX1 fir_data_reg_24__3_ ( .D(fir_data[131]), .CK(clk), .Q(fir_data[115])
         );
  DFFQX1 fir_data_reg_24__2_ ( .D(fir_data[130]), .CK(clk), .Q(fir_data[114])
         );
  DFFQX1 fir_data_reg_24__1_ ( .D(fir_data[129]), .CK(clk), .Q(fir_data[113])
         );
  DFFQX1 fir_data_reg_25__3_ ( .D(fir_data[115]), .CK(clk), .Q(fir_data[99])
         );
  DFFQX1 fir_data_reg_25__2_ ( .D(fir_data[114]), .CK(clk), .Q(fir_data[98])
         );
  DFFQX1 fir_data_reg_25__1_ ( .D(fir_data[113]), .CK(clk), .Q(fir_data[97])
         );
  DFFQX1 fir_data_reg_26__3_ ( .D(fir_data[99]), .CK(clk), .Q(fir_data[83]) );
  DFFQX1 fir_data_reg_26__2_ ( .D(fir_data[98]), .CK(clk), .Q(fir_data[82]) );
  DFFQX1 fir_data_reg_26__1_ ( .D(fir_data[97]), .CK(clk), .Q(fir_data[81]) );
  DFFQX1 fir_data_reg_27__3_ ( .D(fir_data[83]), .CK(clk), .Q(fir_data[67]) );
  DFFQX1 fir_data_reg_27__2_ ( .D(fir_data[82]), .CK(clk), .Q(fir_data[66]) );
  DFFQX1 fir_data_reg_27__1_ ( .D(fir_data[81]), .CK(clk), .Q(fir_data[65]) );
  DFFQX1 fir_data_reg_28__3_ ( .D(fir_data[67]), .CK(clk), .Q(fir_data[51]) );
  DFFQX1 fir_data_reg_28__2_ ( .D(fir_data[66]), .CK(clk), .Q(fir_data[50]) );
  DFFQX1 fir_data_reg_28__1_ ( .D(fir_data[65]), .CK(clk), .Q(fir_data[49]) );
  DFFQX1 fir_data_reg_29__3_ ( .D(fir_data[51]), .CK(clk), .Q(fir_data[35]) );
  DFFQX1 fir_data_reg_29__2_ ( .D(fir_data[50]), .CK(clk), .Q(fir_data[34]) );
  DFFQX1 fir_data_reg_29__1_ ( .D(fir_data[49]), .CK(clk), .Q(fir_data[33]) );
  DFFQX1 fir_data_reg_30__3_ ( .D(fir_data[35]), .CK(clk), .Q(fir_data[19]) );
  DFFQX1 fir_data_reg_30__2_ ( .D(fir_data[34]), .CK(clk), .Q(fir_data[18]) );
  DFFQX1 fir_data_reg_30__1_ ( .D(fir_data[33]), .CK(clk), .Q(fir_data[17]) );
  DFFQX1 fir_data_reg_1__0_ ( .D(fir_data[496]), .CK(clk), .Q(fir_data[480])
         );
  DFFQX1 fir_data_reg_2__0_ ( .D(fir_data[480]), .CK(clk), .Q(fir_data[464])
         );
  DFFQX1 fir_data_reg_3__0_ ( .D(fir_data[464]), .CK(clk), .Q(fir_data[448])
         );
  DFFQX1 fir_data_reg_4__0_ ( .D(fir_data[448]), .CK(clk), .Q(fir_data[432])
         );
  DFFQX1 fir_data_reg_5__0_ ( .D(fir_data[432]), .CK(clk), .Q(fir_data[416])
         );
  DFFQX1 fir_data_reg_6__0_ ( .D(fir_data[416]), .CK(clk), .Q(fir_data[400])
         );
  DFFQX1 fir_data_reg_7__0_ ( .D(fir_data[400]), .CK(clk), .Q(fir_data[384])
         );
  DFFQX1 fir_data_reg_8__0_ ( .D(fir_data[384]), .CK(clk), .Q(fir_data[368])
         );
  DFFQX1 fir_data_reg_9__0_ ( .D(fir_data[368]), .CK(clk), .Q(fir_data[352])
         );
  DFFQX1 fir_data_reg_10__0_ ( .D(fir_data[352]), .CK(clk), .Q(fir_data[336])
         );
  DFFQX1 fir_data_reg_11__0_ ( .D(fir_data[336]), .CK(clk), .Q(fir_data[320])
         );
  DFFQX1 fir_data_reg_12__0_ ( .D(fir_data[320]), .CK(clk), .Q(fir_data[304])
         );
  DFFQX1 fir_data_reg_13__0_ ( .D(fir_data[304]), .CK(clk), .Q(fir_data[288])
         );
  DFFQX1 fir_data_reg_14__0_ ( .D(fir_data[288]), .CK(clk), .Q(fir_data[272])
         );
  DFFQX1 fir_data_reg_15__0_ ( .D(fir_data[272]), .CK(clk), .Q(fir_data[256])
         );
  DFFTRX1 fir_data_reg_0__0_ ( .D(data[0]), .RN(n56), .CK(clk), .Q(
        fir_data[496]) );
  DFFQX1 temp_mul_add_fir_reg_0__20_ ( .D(mul_add_fir[476]), .CK(clk), .Q(
        temp_mul_add_fir[500]) );
  DFFQX1 temp_mul_add_fir_reg_0__19_ ( .D(mul_add_fir[475]), .CK(clk), .Q(
        temp_mul_add_fir[499]) );
  DFFQX1 temp_mul_add_fir_reg_0__18_ ( .D(mul_add_fir[474]), .CK(clk), .Q(
        temp_mul_add_fir[498]) );
  DFFQX1 temp_mul_add_fir_reg_0__17_ ( .D(mul_add_fir[473]), .CK(clk), .Q(
        temp_mul_add_fir[497]) );
  DFFQX1 temp_mul_add_fir_reg_0__16_ ( .D(mul_add_fir[472]), .CK(clk), .Q(
        temp_mul_add_fir[496]) );
  DFFQX1 temp_mul_add_fir_reg_0__15_ ( .D(mul_add_fir[471]), .CK(clk), .Q(
        temp_mul_add_fir[495]) );
  DFFQX1 temp_mul_add_fir_reg_0__14_ ( .D(mul_add_fir[470]), .CK(clk), .Q(
        temp_mul_add_fir[494]) );
  DFFQX1 temp_mul_add_fir_reg_2__19_ ( .D(mul_add_fir[413]), .CK(clk), .Q(
        temp_mul_add_fir[435]) );
  DFFQX1 temp_mul_add_fir_reg_2__18_ ( .D(mul_add_fir[412]), .CK(clk), .Q(
        temp_mul_add_fir[434]) );
  DFFQX1 temp_mul_add_fir_reg_2__17_ ( .D(mul_add_fir[411]), .CK(clk), .Q(
        temp_mul_add_fir[433]) );
  DFFQX1 temp_mul_add_fir_reg_2__16_ ( .D(mul_add_fir[410]), .CK(clk), .Q(
        temp_mul_add_fir[432]) );
  DFFQX1 temp_mul_add_fir_reg_2__15_ ( .D(mul_add_fir[409]), .CK(clk), .Q(
        temp_mul_add_fir[431]) );
  DFFQX1 temp_mul_add_fir_reg_2__14_ ( .D(mul_add_fir[408]), .CK(clk), .Q(
        temp_mul_add_fir[430]) );
  DFFQX1 temp_mul_add_fir_reg_4__19_ ( .D(mul_add_fir[349]), .CK(clk), .Q(
        temp_mul_add_fir[371]) );
  DFFQX1 temp_mul_add_fir_reg_4__18_ ( .D(mul_add_fir[348]), .CK(clk), .Q(
        temp_mul_add_fir[370]) );
  DFFQX1 temp_mul_add_fir_reg_4__17_ ( .D(mul_add_fir[347]), .CK(clk), .Q(
        temp_mul_add_fir[369]) );
  DFFQX1 temp_mul_add_fir_reg_4__16_ ( .D(mul_add_fir[346]), .CK(clk), .Q(
        temp_mul_add_fir[368]) );
  DFFQX1 temp_mul_add_fir_reg_4__15_ ( .D(mul_add_fir[345]), .CK(clk), .Q(
        temp_mul_add_fir[367]) );
  DFFQX1 temp_mul_add_fir_reg_4__14_ ( .D(mul_add_fir[344]), .CK(clk), .Q(
        temp_mul_add_fir[366]) );
  DFFQX1 temp_mul_add_fir_reg_6__19_ ( .D(mul_add_fir[286]), .CK(clk), .Q(
        temp_mul_add_fir[307]) );
  DFFQX1 temp_mul_add_fir_reg_6__18_ ( .D(mul_add_fir[285]), .CK(clk), .Q(
        temp_mul_add_fir[306]) );
  DFFQX1 temp_mul_add_fir_reg_6__17_ ( .D(mul_add_fir[284]), .CK(clk), .Q(
        temp_mul_add_fir[305]) );
  DFFQX1 temp_mul_add_fir_reg_6__16_ ( .D(mul_add_fir[283]), .CK(clk), .Q(
        temp_mul_add_fir[304]) );
  DFFQX1 temp_mul_add_fir_reg_6__15_ ( .D(mul_add_fir[282]), .CK(clk), .Q(
        temp_mul_add_fir[303]) );
  DFFQX1 temp_mul_add_fir_reg_6__14_ ( .D(mul_add_fir[281]), .CK(clk), .Q(
        temp_mul_add_fir[302]) );
  DFFQX1 temp_mul_add_fir_reg_8__19_ ( .D(mul_add_fir[235]), .CK(clk), .Q(
        temp_mul_add_fir[243]) );
  DFFQX1 temp_mul_add_fir_reg_8__18_ ( .D(mul_add_fir[234]), .CK(clk), .Q(
        temp_mul_add_fir[242]) );
  DFFQX1 temp_mul_add_fir_reg_8__17_ ( .D(mul_add_fir[233]), .CK(clk), .Q(
        temp_mul_add_fir[241]) );
  DFFQX1 temp_mul_add_fir_reg_8__16_ ( .D(mul_add_fir[232]), .CK(clk), .Q(
        temp_mul_add_fir[240]) );
  DFFQX1 temp_mul_add_fir_reg_8__15_ ( .D(mul_add_fir[231]), .CK(clk), .Q(
        temp_mul_add_fir[239]) );
  DFFQX1 temp_mul_add_fir_reg_8__14_ ( .D(mul_add_fir[230]), .CK(clk), .Q(
        temp_mul_add_fir[238]) );
  DFFQX1 temp_mul_add_fir_reg_10__19_ ( .D(mul_add_fir[172]), .CK(clk), .Q(
        temp_mul_add_fir[179]) );
  DFFQX1 temp_mul_add_fir_reg_10__18_ ( .D(mul_add_fir[171]), .CK(clk), .Q(
        temp_mul_add_fir[178]) );
  DFFQX1 temp_mul_add_fir_reg_10__17_ ( .D(mul_add_fir[170]), .CK(clk), .Q(
        temp_mul_add_fir[177]) );
  DFFQX1 temp_mul_add_fir_reg_10__16_ ( .D(mul_add_fir[169]), .CK(clk), .Q(
        temp_mul_add_fir[176]) );
  DFFQX1 temp_mul_add_fir_reg_10__15_ ( .D(mul_add_fir[168]), .CK(clk), .Q(
        temp_mul_add_fir[175]) );
  DFFQX1 temp_mul_add_fir_reg_10__14_ ( .D(mul_add_fir[167]), .CK(clk), .Q(
        temp_mul_add_fir[174]) );
  DFFQX1 temp_mul_add_fir_reg_12__19_ ( .D(mul_add_fir[111]), .CK(clk), .Q(
        temp_mul_add_fir[115]) );
  DFFQX1 temp_mul_add_fir_reg_12__18_ ( .D(mul_add_fir[110]), .CK(clk), .Q(
        temp_mul_add_fir[114]) );
  DFFQX1 temp_mul_add_fir_reg_12__17_ ( .D(mul_add_fir[109]), .CK(clk), .Q(
        temp_mul_add_fir[113]) );
  DFFQX1 temp_mul_add_fir_reg_12__16_ ( .D(mul_add_fir[108]), .CK(clk), .Q(
        temp_mul_add_fir[112]) );
  DFFQX1 temp_mul_add_fir_reg_12__15_ ( .D(mul_add_fir[107]), .CK(clk), .Q(
        temp_mul_add_fir[111]) );
  DFFQX1 temp_mul_add_fir_reg_12__14_ ( .D(mul_add_fir[106]), .CK(clk), .Q(
        temp_mul_add_fir[110]) );
  DFFQX1 temp_mul_add_fir_reg_14__19_ ( .D(mul_add_fir[50]), .CK(clk), .Q(
        temp_mul_add_fir[51]) );
  DFFQX1 temp_mul_add_fir_reg_14__18_ ( .D(mul_add_fir[49]), .CK(clk), .Q(
        temp_mul_add_fir[50]) );
  DFFQX1 temp_mul_add_fir_reg_14__17_ ( .D(mul_add_fir[48]), .CK(clk), .Q(
        temp_mul_add_fir[49]) );
  DFFQX1 temp_mul_add_fir_reg_14__16_ ( .D(mul_add_fir[47]), .CK(clk), .Q(
        temp_mul_add_fir[48]) );
  DFFQX1 temp_mul_add_fir_reg_14__15_ ( .D(mul_add_fir[46]), .CK(clk), .Q(
        temp_mul_add_fir[47]) );
  DFFQX1 temp_mul_add_fir_reg_14__14_ ( .D(mul_add_fir[45]), .CK(clk), .Q(
        temp_mul_add_fir[46]) );
  DFFQX1 temp_add_fir_reg_5__15_ ( .D(add_fir[175]), .CK(clk), .Q(
        temp_add_fir[172]) );
  DFFQX1 temp_add_fir_reg_6__15_ ( .D(add_fir[159]), .CK(clk), .Q(
        temp_add_fir[156]) );
  DFFQX1 temp_add_fir_reg_7__11_ ( .D(add_fir[139]), .CK(clk), .Q(
        temp_add_fir[136]) );
  DFFQX1 temp_add_fir_reg_7__10_ ( .D(add_fir[138]), .CK(clk), .Q(
        temp_add_fir[135]) );
  DFFQX1 temp_add_fir_reg_7__9_ ( .D(add_fir[137]), .CK(clk), .Q(
        temp_add_fir[134]) );
  DFFQX1 temp_add_fir_reg_6__14_ ( .D(add_fir[158]), .CK(clk), .Q(
        temp_add_fir[155]) );
  DFFQX1 temp_mul_add_fir_reg_1__19_ ( .D(mul_add_fir[444]), .CK(clk), .Q(
        temp_mul_add_fir[467]) );
  DFFQX1 temp_mul_add_fir_reg_1__18_ ( .D(mul_add_fir[443]), .CK(clk), .Q(
        temp_mul_add_fir[466]) );
  DFFQX1 temp_mul_add_fir_reg_1__17_ ( .D(mul_add_fir[442]), .CK(clk), .Q(
        temp_mul_add_fir[465]) );
  DFFQX1 temp_mul_add_fir_reg_1__16_ ( .D(mul_add_fir[441]), .CK(clk), .Q(
        temp_mul_add_fir[464]) );
  DFFQX1 temp_mul_add_fir_reg_1__15_ ( .D(mul_add_fir[440]), .CK(clk), .Q(
        temp_mul_add_fir[463]) );
  DFFQX1 temp_mul_add_fir_reg_1__14_ ( .D(mul_add_fir[439]), .CK(clk), .Q(
        temp_mul_add_fir[462]) );
  DFFQX1 temp_mul_add_fir_reg_3__19_ ( .D(mul_add_fir[381]), .CK(clk), .Q(
        temp_mul_add_fir[403]) );
  DFFQX1 temp_mul_add_fir_reg_3__18_ ( .D(mul_add_fir[380]), .CK(clk), .Q(
        temp_mul_add_fir[402]) );
  DFFQX1 temp_mul_add_fir_reg_3__17_ ( .D(mul_add_fir[379]), .CK(clk), .Q(
        temp_mul_add_fir[401]) );
  DFFQX1 temp_mul_add_fir_reg_3__16_ ( .D(mul_add_fir[378]), .CK(clk), .Q(
        temp_mul_add_fir[400]) );
  DFFQX1 temp_mul_add_fir_reg_3__15_ ( .D(mul_add_fir[377]), .CK(clk), .Q(
        temp_mul_add_fir[399]) );
  DFFQX1 temp_mul_add_fir_reg_3__14_ ( .D(mul_add_fir[376]), .CK(clk), .Q(
        temp_mul_add_fir[398]) );
  DFFQX1 temp_mul_add_fir_reg_5__19_ ( .D(mul_add_fir[317]), .CK(clk), .Q(
        temp_mul_add_fir[339]) );
  DFFQX1 temp_mul_add_fir_reg_5__18_ ( .D(mul_add_fir[316]), .CK(clk), .Q(
        temp_mul_add_fir[338]) );
  DFFQX1 temp_mul_add_fir_reg_5__17_ ( .D(mul_add_fir[315]), .CK(clk), .Q(
        temp_mul_add_fir[337]) );
  DFFQX1 temp_mul_add_fir_reg_5__16_ ( .D(mul_add_fir[314]), .CK(clk), .Q(
        temp_mul_add_fir[336]) );
  DFFQX1 temp_mul_add_fir_reg_5__15_ ( .D(mul_add_fir[313]), .CK(clk), .Q(
        temp_mul_add_fir[335]) );
  DFFQX1 temp_mul_add_fir_reg_5__14_ ( .D(mul_add_fir[312]), .CK(clk), .Q(
        temp_mul_add_fir[334]) );
  DFFQX1 temp_mul_add_fir_reg_7__19_ ( .D(mul_add_fir[265]), .CK(clk), .Q(
        temp_mul_add_fir[275]) );
  DFFQX1 temp_mul_add_fir_reg_7__18_ ( .D(mul_add_fir[264]), .CK(clk), .Q(
        temp_mul_add_fir[274]) );
  DFFQX1 temp_mul_add_fir_reg_7__17_ ( .D(mul_add_fir[263]), .CK(clk), .Q(
        temp_mul_add_fir[273]) );
  DFFQX1 temp_mul_add_fir_reg_7__16_ ( .D(mul_add_fir[262]), .CK(clk), .Q(
        temp_mul_add_fir[272]) );
  DFFQX1 temp_mul_add_fir_reg_7__15_ ( .D(mul_add_fir[261]), .CK(clk), .Q(
        temp_mul_add_fir[271]) );
  DFFQX1 temp_mul_add_fir_reg_7__14_ ( .D(mul_add_fir[260]), .CK(clk), .Q(
        temp_mul_add_fir[270]) );
  DFFQX1 temp_mul_add_fir_reg_9__19_ ( .D(mul_add_fir[203]), .CK(clk), .Q(
        temp_mul_add_fir[211]) );
  DFFQX1 temp_mul_add_fir_reg_9__18_ ( .D(mul_add_fir[202]), .CK(clk), .Q(
        temp_mul_add_fir[210]) );
  DFFQX1 temp_mul_add_fir_reg_9__17_ ( .D(mul_add_fir[201]), .CK(clk), .Q(
        temp_mul_add_fir[209]) );
  DFFQX1 temp_mul_add_fir_reg_9__16_ ( .D(mul_add_fir[200]), .CK(clk), .Q(
        temp_mul_add_fir[208]) );
  DFFQX1 temp_mul_add_fir_reg_9__15_ ( .D(mul_add_fir[199]), .CK(clk), .Q(
        temp_mul_add_fir[207]) );
  DFFQX1 temp_mul_add_fir_reg_9__14_ ( .D(mul_add_fir[198]), .CK(clk), .Q(
        temp_mul_add_fir[206]) );
  DFFQX1 temp_mul_add_fir_reg_11__19_ ( .D(mul_add_fir[141]), .CK(clk), .Q(
        temp_mul_add_fir[147]) );
  DFFQX1 temp_mul_add_fir_reg_11__18_ ( .D(mul_add_fir[140]), .CK(clk), .Q(
        temp_mul_add_fir[146]) );
  DFFQX1 temp_mul_add_fir_reg_11__17_ ( .D(mul_add_fir[139]), .CK(clk), .Q(
        temp_mul_add_fir[145]) );
  DFFQX1 temp_mul_add_fir_reg_11__16_ ( .D(mul_add_fir[138]), .CK(clk), .Q(
        temp_mul_add_fir[144]) );
  DFFQX1 temp_mul_add_fir_reg_11__15_ ( .D(mul_add_fir[137]), .CK(clk), .Q(
        temp_mul_add_fir[143]) );
  DFFQX1 temp_mul_add_fir_reg_11__14_ ( .D(mul_add_fir[136]), .CK(clk), .Q(
        temp_mul_add_fir[142]) );
  DFFQX1 temp_mul_add_fir_reg_13__19_ ( .D(mul_add_fir[80]), .CK(clk), .Q(
        temp_mul_add_fir[83]) );
  DFFQX1 temp_mul_add_fir_reg_13__18_ ( .D(mul_add_fir[79]), .CK(clk), .Q(
        temp_mul_add_fir[82]) );
  DFFQX1 temp_mul_add_fir_reg_13__17_ ( .D(mul_add_fir[78]), .CK(clk), .Q(
        temp_mul_add_fir[81]) );
  DFFQX1 temp_mul_add_fir_reg_13__16_ ( .D(mul_add_fir[77]), .CK(clk), .Q(
        temp_mul_add_fir[80]) );
  DFFQX1 temp_mul_add_fir_reg_13__15_ ( .D(mul_add_fir[76]), .CK(clk), .Q(
        temp_mul_add_fir[79]) );
  DFFQX1 temp_mul_add_fir_reg_13__14_ ( .D(mul_add_fir[75]), .CK(clk), .Q(
        temp_mul_add_fir[78]) );
  DFFQX1 temp_mul_add_fir_reg_15__19_ ( .D(mul_add_fir[19]), .CK(clk), .Q(
        temp_mul_add_fir[19]) );
  DFFQX1 temp_mul_add_fir_reg_15__18_ ( .D(mul_add_fir[18]), .CK(clk), .Q(
        temp_mul_add_fir[18]) );
  DFFQX1 temp_mul_add_fir_reg_15__17_ ( .D(mul_add_fir[17]), .CK(clk), .Q(
        temp_mul_add_fir[17]) );
  DFFQX1 temp_mul_add_fir_reg_15__16_ ( .D(mul_add_fir[16]), .CK(clk), .Q(
        temp_mul_add_fir[16]) );
  DFFQX1 temp_mul_add_fir_reg_15__15_ ( .D(mul_add_fir[15]), .CK(clk), .Q(
        temp_mul_add_fir[15]) );
  DFFQX1 temp_mul_add_fir_reg_15__14_ ( .D(mul_add_fir[14]), .CK(clk), .Q(
        temp_mul_add_fir[14]) );
  DFFQX1 temp_add_fir_reg_0__15_ ( .D(add_fir[255]), .CK(clk), .Q(
        temp_add_fir[252]) );
  DFFQX1 temp_add_fir_reg_1__15_ ( .D(add_fir[239]), .CK(clk), .Q(
        temp_add_fir[236]) );
  DFFQX1 temp_add_fir_reg_3__14_ ( .D(add_fir[206]), .CK(clk), .Q(
        temp_add_fir[203]) );
  DFFQX1 temp_add_fir_reg_0__14_ ( .D(add_fir[254]), .CK(clk), .Q(
        temp_add_fir[251]) );
  DFFQX1 temp_add_fir_reg_3__15_ ( .D(add_fir[207]), .CK(clk), .Q(
        temp_add_fir[204]) );
  DFFQX1 temp_add_fir_reg_2__15_ ( .D(add_fir[223]), .CK(clk), .Q(
        temp_add_fir[220]) );
  DFFQX1 temp_add_fir_reg_5__14_ ( .D(add_fir[174]), .CK(clk), .Q(
        temp_add_fir[171]) );
  DFFQX1 temp_add_fir_reg_1__13_ ( .D(add_fir[237]), .CK(clk), .Q(
        temp_add_fir[234]) );
  DFFQX1 temp_add_fir_reg_1__14_ ( .D(add_fir[238]), .CK(clk), .Q(
        temp_add_fir[235]) );
  DFFQX1 temp_add_fir_reg_4__14_ ( .D(add_fir[190]), .CK(clk), .Q(
        temp_add_fir[187]) );
  DFFQX1 temp_mul_add_fir_reg_0__13_ ( .D(mul_add_fir[469]), .CK(clk), .Q(
        temp_mul_add_fir[493]) );
  DFFQX1 temp_mul_add_fir_reg_0__12_ ( .D(mul_add_fir[468]), .CK(clk), .Q(
        temp_mul_add_fir[492]) );
  DFFQX1 temp_mul_add_fir_reg_2__13_ ( .D(mul_add_fir[407]), .CK(clk), .Q(
        temp_mul_add_fir[429]) );
  DFFQX1 temp_mul_add_fir_reg_2__12_ ( .D(mul_add_fir[406]), .CK(clk), .Q(
        temp_mul_add_fir[428]) );
  DFFQX1 temp_mul_add_fir_reg_4__13_ ( .D(mul_add_fir[343]), .CK(clk), .Q(
        temp_mul_add_fir[365]) );
  DFFQX1 temp_mul_add_fir_reg_4__12_ ( .D(mul_add_fir[342]), .CK(clk), .Q(
        temp_mul_add_fir[364]) );
  DFFQX1 temp_mul_add_fir_reg_6__13_ ( .D(mul_add_fir[280]), .CK(clk), .Q(
        temp_mul_add_fir[301]) );
  DFFQX1 temp_mul_add_fir_reg_6__12_ ( .D(mul_add_fir[279]), .CK(clk), .Q(
        temp_mul_add_fir[300]) );
  DFFQX1 temp_mul_add_fir_reg_8__13_ ( .D(mul_add_fir[229]), .CK(clk), .Q(
        temp_mul_add_fir[237]) );
  DFFQX1 temp_mul_add_fir_reg_8__12_ ( .D(mul_add_fir[228]), .CK(clk), .Q(
        temp_mul_add_fir[236]) );
  DFFQX1 temp_mul_add_fir_reg_10__13_ ( .D(mul_add_fir[166]), .CK(clk), .Q(
        temp_mul_add_fir[173]) );
  DFFQX1 temp_mul_add_fir_reg_10__12_ ( .D(mul_add_fir[165]), .CK(clk), .Q(
        temp_mul_add_fir[172]) );
  DFFQX1 temp_mul_add_fir_reg_12__13_ ( .D(mul_add_fir[105]), .CK(clk), .Q(
        temp_mul_add_fir[109]) );
  DFFQX1 temp_mul_add_fir_reg_12__12_ ( .D(mul_add_fir[104]), .CK(clk), .Q(
        temp_mul_add_fir[108]) );
  DFFQX1 temp_mul_add_fir_reg_14__13_ ( .D(mul_add_fir[44]), .CK(clk), .Q(
        temp_mul_add_fir[45]) );
  DFFQX1 temp_mul_add_fir_reg_14__12_ ( .D(mul_add_fir[43]), .CK(clk), .Q(
        temp_mul_add_fir[44]) );
  DFFQX1 temp_add_fir_reg_4__15_ ( .D(add_fir[191]), .CK(clk), .Q(
        temp_add_fir[188]) );
  DFFQX1 temp_add_fir_reg_12__15_ ( .D(add_fir[63]), .CK(clk), .Q(
        temp_add_fir[63]) );
  DFFQX1 temp_add_fir_reg_3__11_ ( .D(add_fir[203]), .CK(clk), .Q(
        temp_add_fir[200]) );
  DFFQX1 temp_add_fir_reg_7__8_ ( .D(add_fir[136]), .CK(clk), .Q(
        temp_add_fir[133]) );
  DFFQX1 temp_add_fir_reg_7__7_ ( .D(add_fir[135]), .CK(clk), .Q(
        temp_add_fir[132]) );
  DFFQX1 temp_add_fir_reg_7__6_ ( .D(add_fir[134]), .CK(clk), .Q(
        temp_add_fir[131]) );
  DFFQX1 temp_add_fir_reg_3__12_ ( .D(add_fir[204]), .CK(clk), .Q(
        temp_add_fir[201]) );
  DFFQX1 temp_add_fir_reg_0__13_ ( .D(add_fir[253]), .CK(clk), .Q(
        temp_add_fir[250]) );
  DFFQX1 temp_add_fir_reg_11__12_ ( .D(add_fir[76]), .CK(clk), .Q(
        temp_add_fir[76]) );
  DFFQX1 temp_add_fir_reg_6__13_ ( .D(add_fir[157]), .CK(clk), .Q(
        temp_add_fir[154]) );
  DFFQX1 temp_add_fir_reg_6__12_ ( .D(add_fir[156]), .CK(clk), .Q(
        temp_add_fir[153]) );
  DFFQX1 temp_add_fir_reg_6__11_ ( .D(add_fir[155]), .CK(clk), .Q(
        temp_add_fir[152]) );
  DFFQX1 temp_mul_add_fir_reg_1__13_ ( .D(mul_add_fir[438]), .CK(clk), .Q(
        temp_mul_add_fir[461]) );
  DFFQX1 temp_mul_add_fir_reg_1__12_ ( .D(mul_add_fir[437]), .CK(clk), .Q(
        temp_mul_add_fir[460]) );
  DFFQX1 temp_mul_add_fir_reg_3__13_ ( .D(mul_add_fir[375]), .CK(clk), .Q(
        temp_mul_add_fir[397]) );
  DFFQX1 temp_mul_add_fir_reg_3__12_ ( .D(mul_add_fir[374]), .CK(clk), .Q(
        temp_mul_add_fir[396]) );
  DFFQX1 temp_mul_add_fir_reg_5__13_ ( .D(mul_add_fir[311]), .CK(clk), .Q(
        temp_mul_add_fir[333]) );
  DFFQX1 temp_mul_add_fir_reg_5__12_ ( .D(mul_add_fir[310]), .CK(clk), .Q(
        temp_mul_add_fir[332]) );
  DFFQX1 temp_mul_add_fir_reg_7__13_ ( .D(mul_add_fir[259]), .CK(clk), .Q(
        temp_mul_add_fir[269]) );
  DFFQX1 temp_mul_add_fir_reg_7__12_ ( .D(mul_add_fir[258]), .CK(clk), .Q(
        temp_mul_add_fir[268]) );
  DFFQX1 temp_mul_add_fir_reg_9__13_ ( .D(mul_add_fir[197]), .CK(clk), .Q(
        temp_mul_add_fir[205]) );
  DFFQX1 temp_mul_add_fir_reg_9__12_ ( .D(mul_add_fir[196]), .CK(clk), .Q(
        temp_mul_add_fir[204]) );
  DFFQX1 temp_mul_add_fir_reg_11__13_ ( .D(mul_add_fir[135]), .CK(clk), .Q(
        temp_mul_add_fir[141]) );
  DFFQX1 temp_mul_add_fir_reg_11__12_ ( .D(mul_add_fir[134]), .CK(clk), .Q(
        temp_mul_add_fir[140]) );
  DFFQX1 temp_mul_add_fir_reg_13__13_ ( .D(mul_add_fir[74]), .CK(clk), .Q(
        temp_mul_add_fir[77]) );
  DFFQX1 temp_mul_add_fir_reg_13__12_ ( .D(mul_add_fir[73]), .CK(clk), .Q(
        temp_mul_add_fir[76]) );
  DFFQX1 temp_mul_add_fir_reg_15__13_ ( .D(mul_add_fir[13]), .CK(clk), .Q(
        temp_mul_add_fir[13]) );
  DFFQX1 temp_mul_add_fir_reg_15__12_ ( .D(mul_add_fir[12]), .CK(clk), .Q(
        temp_mul_add_fir[12]) );
  DFFQX1 temp_add_fir_reg_3__13_ ( .D(add_fir[205]), .CK(clk), .Q(
        temp_add_fir[202]) );
  DFFQX1 temp_add_fir_reg_1__10_ ( .D(add_fir[234]), .CK(clk), .Q(
        temp_add_fir[231]) );
  DFFQX1 temp_add_fir_reg_0__12_ ( .D(add_fir[252]), .CK(clk), .Q(
        temp_add_fir[249]) );
  DFFQX1 temp_add_fir_reg_0__11_ ( .D(add_fir[251]), .CK(clk), .Q(
        temp_add_fir[248]) );
  DFFQX1 temp_add_fir_reg_11__13_ ( .D(add_fir[77]), .CK(clk), .Q(
        temp_add_fir[77]) );
  DFFQX1 temp_add_fir_reg_2__13_ ( .D(add_fir[221]), .CK(clk), .Q(
        temp_add_fir[218]) );
  DFFQX1 temp_add_fir_reg_5__12_ ( .D(add_fir[172]), .CK(clk), .Q(
        temp_add_fir[169]) );
  DFFQX1 temp_add_fir_reg_5__13_ ( .D(add_fir[173]), .CK(clk), .Q(
        temp_add_fir[170]) );
  DFFQX1 temp_add_fir_reg_1__12_ ( .D(add_fir[236]), .CK(clk), .Q(
        temp_add_fir[233]) );
  DFFQX1 temp_add_fir_reg_1__11_ ( .D(add_fir[235]), .CK(clk), .Q(
        temp_add_fir[232]) );
  DFFQX1 temp_add_fir_reg_5__11_ ( .D(add_fir[171]), .CK(clk), .Q(
        temp_add_fir[168]) );
  DFFQX1 temp_add_fir_reg_5__10_ ( .D(add_fir[170]), .CK(clk), .Q(
        temp_add_fir[167]) );
  DFFQX1 temp_add_fir_reg_2__14_ ( .D(add_fir[222]), .CK(clk), .Q(
        temp_add_fir[219]) );
  DFFQX1 temp_add_fir_reg_10__15_ ( .D(add_fir[95]), .CK(clk), .Q(
        temp_add_fir[95]) );
  DFFQX1 temp_add_fir_reg_2__12_ ( .D(add_fir[220]), .CK(clk), .Q(
        temp_add_fir[217]) );
  DFFQX1 temp_add_fir_reg_4__13_ ( .D(add_fir[189]), .CK(clk), .Q(
        temp_add_fir[186]) );
  DFFQX1 temp_add_fir_reg_4__11_ ( .D(add_fir[187]), .CK(clk), .Q(
        temp_add_fir[184]) );
  DFFQX1 temp_add_fir_reg_11__14_ ( .D(add_fir[78]), .CK(clk), .Q(
        temp_add_fir[78]) );
  DFFQX1 temp_add_fir_reg_4__12_ ( .D(add_fir[188]), .CK(clk), .Q(
        temp_add_fir[185]) );
  DFFQX1 temp_add_fir_reg_11__15_ ( .D(add_fir[79]), .CK(clk), .Q(
        temp_add_fir[79]) );
  DFFQX1 temp_add_fir_reg_12__14_ ( .D(add_fir[62]), .CK(clk), .Q(
        temp_add_fir[62]) );
  DFFQX1 temp_mul_add_fir_reg_0__11_ ( .D(mul_add_fir[467]), .CK(clk), .Q(
        temp_mul_add_fir[491]) );
  DFFQX1 temp_mul_add_fir_reg_0__10_ ( .D(mul_add_fir[466]), .CK(clk), .Q(
        temp_mul_add_fir[490]) );
  DFFQX1 temp_mul_add_fir_reg_2__11_ ( .D(mul_add_fir[405]), .CK(clk), .Q(
        temp_mul_add_fir[427]) );
  DFFQX1 temp_mul_add_fir_reg_2__10_ ( .D(mul_add_fir[404]), .CK(clk), .Q(
        temp_mul_add_fir[426]) );
  DFFQX1 temp_mul_add_fir_reg_4__11_ ( .D(mul_add_fir[341]), .CK(clk), .Q(
        temp_mul_add_fir[363]) );
  DFFQX1 temp_mul_add_fir_reg_4__10_ ( .D(mul_add_fir[340]), .CK(clk), .Q(
        temp_mul_add_fir[362]) );
  DFFQX1 temp_mul_add_fir_reg_6__11_ ( .D(mul_add_fir[278]), .CK(clk), .Q(
        temp_mul_add_fir[299]) );
  DFFQX1 temp_mul_add_fir_reg_6__10_ ( .D(mul_add_fir[277]), .CK(clk), .Q(
        temp_mul_add_fir[298]) );
  DFFQX1 temp_mul_add_fir_reg_8__11_ ( .D(mul_add_fir[227]), .CK(clk), .Q(
        temp_mul_add_fir[235]) );
  DFFQX1 temp_mul_add_fir_reg_8__10_ ( .D(mul_add_fir[226]), .CK(clk), .Q(
        temp_mul_add_fir[234]) );
  DFFQX1 temp_mul_add_fir_reg_8__9_ ( .D(mul_add_fir[225]), .CK(clk), .Q(
        temp_mul_add_fir[233]) );
  DFFQX1 temp_mul_add_fir_reg_10__11_ ( .D(mul_add_fir[164]), .CK(clk), .Q(
        temp_mul_add_fir[171]) );
  DFFQX1 temp_mul_add_fir_reg_10__10_ ( .D(mul_add_fir[163]), .CK(clk), .Q(
        temp_mul_add_fir[170]) );
  DFFQX1 temp_mul_add_fir_reg_10__9_ ( .D(mul_add_fir[162]), .CK(clk), .Q(
        temp_mul_add_fir[169]) );
  DFFQX1 temp_mul_add_fir_reg_12__11_ ( .D(mul_add_fir[103]), .CK(clk), .Q(
        temp_mul_add_fir[107]) );
  DFFQX1 temp_mul_add_fir_reg_12__10_ ( .D(mul_add_fir[102]), .CK(clk), .Q(
        temp_mul_add_fir[106]) );
  DFFQX1 temp_mul_add_fir_reg_12__9_ ( .D(mul_add_fir[101]), .CK(clk), .Q(
        temp_mul_add_fir[105]) );
  DFFQX1 temp_mul_add_fir_reg_14__11_ ( .D(mul_add_fir[42]), .CK(clk), .Q(
        temp_mul_add_fir[43]) );
  DFFQX1 temp_mul_add_fir_reg_14__10_ ( .D(mul_add_fir[41]), .CK(clk), .Q(
        temp_mul_add_fir[42]) );
  DFFQX1 temp_mul_add_fir_reg_14__9_ ( .D(mul_add_fir[40]), .CK(clk), .Q(
        temp_mul_add_fir[41]) );
  DFFQX1 temp_add_fir_reg_3__9_ ( .D(add_fir[201]), .CK(clk), .Q(
        temp_add_fir[198]) );
  DFFQX1 temp_add_fir_reg_7__5_ ( .D(add_fir[133]), .CK(clk), .Q(
        temp_add_fir[130]) );
  DFFQX1 temp_add_fir_reg_7__4_ ( .D(add_fir[132]), .CK(clk), .Q(
        temp_add_fir[129]) );
  DFFQX1 temp_add_fir_reg_7__2_ ( .D(add_fir[130]), .CK(clk), .Q(
        mul_add_fir[250]) );
  DFFQX1 temp_add_fir_reg_7__1_ ( .D(add_fir[129]), .CK(clk), .Q(
        mul_add_fir[249]) );
  DFFQX1 temp_add_fir_reg_7__3_ ( .D(add_fir[131]), .CK(clk), .Q(
        temp_add_fir[128]) );
  DFFQX1 temp_add_fir_reg_0__8_ ( .D(add_fir[248]), .CK(clk), .Q(
        temp_add_fir[245]) );
  DFFQX1 temp_add_fir_reg_3__10_ ( .D(add_fir[202]), .CK(clk), .Q(
        temp_add_fir[199]) );
  DFFQX1 temp_add_fir_reg_3__8_ ( .D(add_fir[200]), .CK(clk), .Q(
        temp_add_fir[197]) );
  DFFQX1 temp_add_fir_reg_11__11_ ( .D(add_fir[75]), .CK(clk), .Q(
        temp_add_fir[75]) );
  DFFQX1 temp_add_fir_reg_11__10_ ( .D(add_fir[74]), .CK(clk), .Q(
        temp_add_fir[74]) );
  DFFQX1 temp_add_fir_reg_11__9_ ( .D(add_fir[73]), .CK(clk), .Q(
        temp_add_fir[73]) );
  DFFQX1 temp_add_fir_reg_6__3_ ( .D(add_fir[147]), .CK(clk), .Q(
        temp_add_fir[144]) );
  DFFQX1 temp_add_fir_reg_6__2_ ( .D(add_fir[146]), .CK(clk), .Q(
        temp_add_fir[143]) );
  DFFQX1 temp_add_fir_reg_6__6_ ( .D(add_fir[150]), .CK(clk), .Q(
        temp_add_fir[147]) );
  DFFQX1 temp_add_fir_reg_7__0_ ( .D(add_fir[128]), .CK(clk), .Q(
        mul_add_fir[248]) );
  DFFQX1 temp_add_fir_reg_6__7_ ( .D(add_fir[151]), .CK(clk), .Q(
        temp_add_fir[148]) );
  DFFQX1 temp_add_fir_reg_6__10_ ( .D(add_fir[154]), .CK(clk), .Q(
        temp_add_fir[151]) );
  DFFQX1 temp_add_fir_reg_6__9_ ( .D(add_fir[153]), .CK(clk), .Q(
        temp_add_fir[150]) );
  DFFQX1 temp_add_fir_reg_6__8_ ( .D(add_fir[152]), .CK(clk), .Q(
        temp_add_fir[149]) );
  DFFQX1 temp_mul_add_fir_reg_1__11_ ( .D(mul_add_fir[436]), .CK(clk), .Q(
        temp_mul_add_fir[459]) );
  DFFQX1 temp_mul_add_fir_reg_1__10_ ( .D(mul_add_fir[435]), .CK(clk), .Q(
        temp_mul_add_fir[458]) );
  DFFQX1 temp_mul_add_fir_reg_3__11_ ( .D(mul_add_fir[373]), .CK(clk), .Q(
        temp_mul_add_fir[395]) );
  DFFQX1 temp_mul_add_fir_reg_3__10_ ( .D(mul_add_fir[372]), .CK(clk), .Q(
        temp_mul_add_fir[394]) );
  DFFQX1 temp_mul_add_fir_reg_5__11_ ( .D(mul_add_fir[309]), .CK(clk), .Q(
        temp_mul_add_fir[331]) );
  DFFQX1 temp_mul_add_fir_reg_5__10_ ( .D(mul_add_fir[308]), .CK(clk), .Q(
        temp_mul_add_fir[330]) );
  DFFQX1 temp_mul_add_fir_reg_7__11_ ( .D(mul_add_fir[257]), .CK(clk), .Q(
        temp_mul_add_fir[267]) );
  DFFQX1 temp_mul_add_fir_reg_7__10_ ( .D(mul_add_fir[256]), .CK(clk), .Q(
        temp_mul_add_fir[266]) );
  DFFQX1 temp_mul_add_fir_reg_9__11_ ( .D(mul_add_fir[195]), .CK(clk), .Q(
        temp_mul_add_fir[203]) );
  DFFQX1 temp_mul_add_fir_reg_9__10_ ( .D(mul_add_fir[194]), .CK(clk), .Q(
        temp_mul_add_fir[202]) );
  DFFQX1 temp_mul_add_fir_reg_9__9_ ( .D(mul_add_fir[193]), .CK(clk), .Q(
        temp_mul_add_fir[201]) );
  DFFQX1 temp_mul_add_fir_reg_11__11_ ( .D(mul_add_fir[133]), .CK(clk), .Q(
        temp_mul_add_fir[139]) );
  DFFQX1 temp_mul_add_fir_reg_11__10_ ( .D(mul_add_fir[132]), .CK(clk), .Q(
        temp_mul_add_fir[138]) );
  DFFQX1 temp_mul_add_fir_reg_11__9_ ( .D(mul_add_fir[131]), .CK(clk), .Q(
        temp_mul_add_fir[137]) );
  DFFQX1 temp_mul_add_fir_reg_13__11_ ( .D(mul_add_fir[72]), .CK(clk), .Q(
        temp_mul_add_fir[75]) );
  DFFQX1 temp_mul_add_fir_reg_13__10_ ( .D(mul_add_fir[71]), .CK(clk), .Q(
        temp_mul_add_fir[74]) );
  DFFQX1 temp_mul_add_fir_reg_13__9_ ( .D(mul_add_fir[70]), .CK(clk), .Q(
        temp_mul_add_fir[73]) );
  DFFQX1 temp_mul_add_fir_reg_15__11_ ( .D(mul_add_fir[11]), .CK(clk), .Q(
        temp_mul_add_fir[11]) );
  DFFQX1 temp_mul_add_fir_reg_15__10_ ( .D(mul_add_fir[10]), .CK(clk), .Q(
        temp_mul_add_fir[10]) );
  DFFQX1 temp_mul_add_fir_reg_15__9_ ( .D(mul_add_fir[9]), .CK(clk), .Q(
        temp_mul_add_fir[9]) );
  DFFQX1 temp_add_fir_reg_1__6_ ( .D(add_fir[230]), .CK(clk), .Q(
        temp_add_fir[227]) );
  DFFQX1 temp_add_fir_reg_1__9_ ( .D(add_fir[233]), .CK(clk), .Q(
        temp_add_fir[230]) );
  DFFQX1 temp_add_fir_reg_1__8_ ( .D(add_fir[232]), .CK(clk), .Q(
        temp_add_fir[229]) );
  DFFQX1 temp_add_fir_reg_1__7_ ( .D(add_fir[231]), .CK(clk), .Q(
        temp_add_fir[228]) );
  DFFQX1 temp_add_fir_reg_0__10_ ( .D(add_fir[250]), .CK(clk), .Q(
        temp_add_fir[247]) );
  DFFQX1 temp_add_fir_reg_0__9_ ( .D(add_fir[249]), .CK(clk), .Q(
        temp_add_fir[246]) );
  DFFQX1 temp_add_fir_reg_0__6_ ( .D(add_fir[246]), .CK(clk), .Q(
        temp_add_fir[243]) );
  DFFQX1 temp_add_fir_reg_2__11_ ( .D(add_fir[219]), .CK(clk), .Q(
        temp_add_fir[216]) );
  DFFQX1 temp_add_fir_reg_14__15_ ( .D(add_fir[31]), .CK(clk), .Q(
        temp_add_fir[31]) );
  DFFQX1 temp_add_fir_reg_5__9_ ( .D(add_fir[169]), .CK(clk), .Q(
        temp_add_fir[166]) );
  DFFQX1 temp_add_fir_reg_5__8_ ( .D(add_fir[168]), .CK(clk), .Q(
        temp_add_fir[165]) );
  DFFQX1 temp_add_fir_reg_8__15_ ( .D(add_fir[127]), .CK(clk), .Q(
        temp_add_fir[127]) );
  DFFQX1 temp_add_fir_reg_9__15_ ( .D(add_fir[111]), .CK(clk), .Q(
        temp_add_fir[111]) );
  DFFQX1 temp_add_fir_reg_9__12_ ( .D(add_fir[108]), .CK(clk), .Q(
        temp_add_fir[108]) );
  DFFQX1 temp_add_fir_reg_10__13_ ( .D(add_fir[93]), .CK(clk), .Q(
        temp_add_fir[93]) );
  DFFQX1 temp_add_fir_reg_2__10_ ( .D(add_fir[218]), .CK(clk), .Q(
        temp_add_fir[215]) );
  DFFQX1 temp_add_fir_reg_2__9_ ( .D(add_fir[217]), .CK(clk), .Q(
        temp_add_fir[214]) );
  DFFQX1 temp_add_fir_reg_4__7_ ( .D(add_fir[183]), .CK(clk), .Q(
        temp_add_fir[180]) );
  DFFQX1 temp_add_fir_reg_8__14_ ( .D(add_fir[126]), .CK(clk), .Q(
        temp_add_fir[126]) );
  DFFQX1 temp_add_fir_reg_8__13_ ( .D(add_fir[125]), .CK(clk), .Q(
        temp_add_fir[125]) );
  DFFQX1 temp_add_fir_reg_9__14_ ( .D(add_fir[110]), .CK(clk), .Q(
        temp_add_fir[110]) );
  DFFQX1 temp_add_fir_reg_9__13_ ( .D(add_fir[109]), .CK(clk), .Q(
        temp_add_fir[109]) );
  DFFQX1 temp_add_fir_reg_8__12_ ( .D(add_fir[124]), .CK(clk), .Q(
        temp_add_fir[124]) );
  DFFQX1 temp_add_fir_reg_4__10_ ( .D(add_fir[186]), .CK(clk), .Q(
        temp_add_fir[183]) );
  DFFQX1 temp_add_fir_reg_4__9_ ( .D(add_fir[185]), .CK(clk), .Q(
        temp_add_fir[182]) );
  DFFQX1 temp_add_fir_reg_4__8_ ( .D(add_fir[184]), .CK(clk), .Q(
        temp_add_fir[181]) );
  DFFQX1 temp_add_fir_reg_10__14_ ( .D(add_fir[94]), .CK(clk), .Q(
        temp_add_fir[94]) );
  DFFQX1 temp_add_fir_reg_13__15_ ( .D(add_fir[47]), .CK(clk), .Q(
        temp_add_fir[47]) );
  DFFQX2 temp_add_fir_reg_12__13_ ( .D(add_fir[61]), .CK(clk), .Q(
        temp_add_fir[61]) );
  DFFQX2 temp_add_fir_reg_12__12_ ( .D(add_fir[60]), .CK(clk), .Q(
        temp_add_fir[60]) );
  DFFQX2 temp_add_fir_reg_12__10_ ( .D(add_fir[58]), .CK(clk), .Q(
        temp_add_fir[58]) );
  DFFQX2 temp_add_fir_reg_12__11_ ( .D(add_fir[59]), .CK(clk), .Q(
        temp_add_fir[59]) );
  DFFQX1 temp_mul_add_fir_reg_0__9_ ( .D(mul_add_fir[465]), .CK(clk), .Q(
        temp_mul_add_fir[489]) );
  DFFQX1 temp_mul_add_fir_reg_0__8_ ( .D(mul_add_fir[464]), .CK(clk), .Q(
        temp_mul_add_fir[488]) );
  DFFQX1 temp_mul_add_fir_reg_2__9_ ( .D(mul_add_fir[403]), .CK(clk), .Q(
        temp_mul_add_fir[425]) );
  DFFQX1 temp_mul_add_fir_reg_4__9_ ( .D(mul_add_fir[339]), .CK(clk), .Q(
        temp_mul_add_fir[361]) );
  DFFQX1 temp_mul_add_fir_reg_4__8_ ( .D(mul_add_fir[338]), .CK(clk), .Q(
        temp_mul_add_fir[360]) );
  DFFQX1 temp_mul_add_fir_reg_6__9_ ( .D(mul_add_fir[276]), .CK(clk), .Q(
        temp_mul_add_fir[297]) );
  DFFQX1 temp_mul_add_fir_reg_8__8_ ( .D(mul_add_fir[224]), .CK(clk), .Q(
        temp_mul_add_fir[232]) );
  DFFQX1 temp_mul_add_fir_reg_12__8_ ( .D(mul_add_fir[100]), .CK(clk), .Q(
        temp_mul_add_fir[104]) );
  DFFQX1 temp_add_fir_reg_0__1_ ( .D(add_fir[241]), .CK(clk), .Q(
        temp_add_fir[238]) );
  DFFQX1 temp_add_fir_reg_11__7_ ( .D(add_fir[71]), .CK(clk), .Q(
        temp_add_fir[71]) );
  DFFQX1 temp_add_fir_reg_11__4_ ( .D(add_fir[68]), .CK(clk), .Q(
        temp_add_fir[68]) );
  DFFQX1 temp_add_fir_reg_13__11_ ( .D(add_fir[43]), .CK(clk), .Q(
        temp_add_fir[43]) );
  DFFQX1 temp_add_fir_reg_0__2_ ( .D(add_fir[242]), .CK(clk), .Q(
        temp_add_fir[239]) );
  DFFQX1 temp_add_fir_reg_11__5_ ( .D(add_fir[69]), .CK(clk), .Q(
        temp_add_fir[69]) );
  DFFQX1 temp_add_fir_reg_13__12_ ( .D(add_fir[44]), .CK(clk), .Q(
        temp_add_fir[44]) );
  DFFQX1 temp_add_fir_reg_0__7_ ( .D(add_fir[247]), .CK(clk), .Q(
        temp_add_fir[244]) );
  DFFQX1 temp_add_fir_reg_0__5_ ( .D(add_fir[245]), .CK(clk), .Q(
        temp_add_fir[242]) );
  DFFQX1 temp_add_fir_reg_0__4_ ( .D(add_fir[244]), .CK(clk), .Q(
        temp_add_fir[241]) );
  DFFQX1 temp_add_fir_reg_0__3_ ( .D(add_fir[243]), .CK(clk), .Q(
        temp_add_fir[240]) );
  DFFQX1 temp_add_fir_reg_3__7_ ( .D(add_fir[199]), .CK(clk), .Q(
        temp_add_fir[196]) );
  DFFQX1 temp_add_fir_reg_3__6_ ( .D(add_fir[198]), .CK(clk), .Q(
        temp_add_fir[195]) );
  DFFQX1 temp_add_fir_reg_3__5_ ( .D(add_fir[197]), .CK(clk), .Q(
        temp_add_fir[194]) );
  DFFQX1 temp_add_fir_reg_3__4_ ( .D(add_fir[196]), .CK(clk), .Q(
        temp_add_fir[193]) );
  DFFQX1 temp_add_fir_reg_3__3_ ( .D(add_fir[195]), .CK(clk), .Q(
        temp_add_fir[192]) );
  DFFQX1 temp_add_fir_reg_11__6_ ( .D(add_fir[70]), .CK(clk), .Q(
        temp_add_fir[70]) );
  DFFQX1 temp_add_fir_reg_13__10_ ( .D(add_fir[42]), .CK(clk), .Q(
        temp_add_fir[42]) );
  DFFQX1 temp_add_fir_reg_11__8_ ( .D(add_fir[72]), .CK(clk), .Q(
        temp_add_fir[72]) );
  DFFQX1 temp_add_fir_reg_6__1_ ( .D(add_fir[145]), .CK(clk), .Q(
        temp_add_fir[142]) );
  DFFQX1 temp_add_fir_reg_6__0_ ( .D(add_fir[144]), .CK(clk), .Q(
        temp_add_fir[141]) );
  DFFQX1 temp_add_fir_reg_6__5_ ( .D(add_fir[149]), .CK(clk), .Q(
        temp_add_fir[146]) );
  DFFQX1 temp_add_fir_reg_6__4_ ( .D(add_fir[148]), .CK(clk), .Q(
        temp_add_fir[145]) );
  DFFQX1 temp_mul_add_fir_reg_1__9_ ( .D(mul_add_fir[434]), .CK(clk), .Q(
        temp_mul_add_fir[457]) );
  DFFQX1 temp_mul_add_fir_reg_1__8_ ( .D(mul_add_fir[433]), .CK(clk), .Q(
        temp_mul_add_fir[456]) );
  DFFQX1 temp_mul_add_fir_reg_3__9_ ( .D(mul_add_fir[371]), .CK(clk), .Q(
        temp_mul_add_fir[393]) );
  DFFQX1 temp_mul_add_fir_reg_5__9_ ( .D(mul_add_fir[307]), .CK(clk), .Q(
        temp_mul_add_fir[329]) );
  DFFQX1 temp_mul_add_fir_reg_7__9_ ( .D(mul_add_fir[255]), .CK(clk), .Q(
        temp_mul_add_fir[265]) );
  DFFQX1 temp_add_fir_reg_1__5_ ( .D(add_fir[229]), .CK(clk), .Q(
        temp_add_fir[226]) );
  DFFQX1 temp_add_fir_reg_1__4_ ( .D(add_fir[228]), .CK(clk), .Q(
        temp_add_fir[225]) );
  DFFQX1 temp_add_fir_reg_1__3_ ( .D(add_fir[227]), .CK(clk), .Q(
        temp_add_fir[224]) );
  DFFQX1 temp_add_fir_reg_8__8_ ( .D(add_fir[120]), .CK(clk), .Q(
        temp_add_fir[120]) );
  DFFQX1 temp_add_fir_reg_9__8_ ( .D(add_fir[104]), .CK(clk), .Q(
        temp_add_fir[104]) );
  DFFQX1 temp_add_fir_reg_10__11_ ( .D(add_fir[91]), .CK(clk), .Q(
        temp_add_fir[91]) );
  DFFQX1 temp_add_fir_reg_15__15_ ( .D(add_fir[15]), .CK(clk), .Q(
        temp_add_fir[15]) );
  DFFQX1 temp_add_fir_reg_2__4_ ( .D(add_fir[212]), .CK(clk), .Q(
        temp_add_fir[209]) );
  DFFQX1 temp_add_fir_reg_9__10_ ( .D(add_fir[106]), .CK(clk), .Q(
        temp_add_fir[106]) );
  DFFQX1 temp_add_fir_reg_14__13_ ( .D(add_fir[29]), .CK(clk), .Q(
        temp_add_fir[29]) );
  DFFQX1 temp_add_fir_reg_5__0_ ( .D(add_fir[160]), .CK(clk), .Q(
        temp_add_fir[157]) );
  DFFQX1 temp_add_fir_reg_8__9_ ( .D(add_fir[121]), .CK(clk), .Q(
        temp_add_fir[121]) );
  DFFQX1 temp_add_fir_reg_9__9_ ( .D(add_fir[105]), .CK(clk), .Q(
        temp_add_fir[105]) );
  DFFQX1 temp_add_fir_reg_2__6_ ( .D(add_fir[214]), .CK(clk), .Q(
        temp_add_fir[211]) );
  DFFQX1 temp_add_fir_reg_2__5_ ( .D(add_fir[213]), .CK(clk), .Q(
        temp_add_fir[210]) );
  DFFQX1 temp_add_fir_reg_8__11_ ( .D(add_fir[123]), .CK(clk), .Q(
        temp_add_fir[123]) );
  DFFQX1 temp_add_fir_reg_5__1_ ( .D(add_fir[161]), .CK(clk), .Q(
        temp_add_fir[158]) );
  DFFQX1 temp_add_fir_reg_5__2_ ( .D(add_fir[162]), .CK(clk), .Q(
        temp_add_fir[159]) );
  DFFQX1 temp_add_fir_reg_5__3_ ( .D(add_fir[163]), .CK(clk), .Q(
        temp_add_fir[160]) );
  DFFQX1 temp_add_fir_reg_13__13_ ( .D(add_fir[45]), .CK(clk), .Q(
        temp_add_fir[45]) );
  DFFQX1 temp_add_fir_reg_10__9_ ( .D(add_fir[89]), .CK(clk), .Q(
        temp_add_fir[89]) );
  DFFQX1 temp_add_fir_reg_5__6_ ( .D(add_fir[166]), .CK(clk), .Q(
        temp_add_fir[163]) );
  DFFQX1 temp_add_fir_reg_5__4_ ( .D(add_fir[164]), .CK(clk), .Q(
        temp_add_fir[161]) );
  DFFQX1 temp_add_fir_reg_5__5_ ( .D(add_fir[165]), .CK(clk), .Q(
        temp_add_fir[162]) );
  DFFQX1 temp_add_fir_reg_5__7_ ( .D(add_fir[167]), .CK(clk), .Q(
        temp_add_fir[164]) );
  DFFQX1 temp_add_fir_reg_14__12_ ( .D(add_fir[28]), .CK(clk), .Q(
        temp_add_fir[28]) );
  DFFQX1 temp_add_fir_reg_14__11_ ( .D(add_fir[27]), .CK(clk), .Q(
        temp_add_fir[27]) );
  DFFQX1 temp_add_fir_reg_2__7_ ( .D(add_fir[215]), .CK(clk), .Q(
        temp_add_fir[212]) );
  DFFQX1 temp_add_fir_reg_4__5_ ( .D(add_fir[181]), .CK(clk), .Q(
        temp_add_fir[178]) );
  DFFQX1 temp_add_fir_reg_4__6_ ( .D(add_fir[182]), .CK(clk), .Q(
        temp_add_fir[179]) );
  DFFQX1 temp_add_fir_reg_8__10_ ( .D(add_fir[122]), .CK(clk), .Q(
        temp_add_fir[122]) );
  DFFQX1 temp_add_fir_reg_14__14_ ( .D(add_fir[30]), .CK(clk), .Q(
        temp_add_fir[30]) );
  DFFQX1 temp_add_fir_reg_2__8_ ( .D(add_fir[216]), .CK(clk), .Q(
        temp_add_fir[213]) );
  DFFQX1 temp_add_fir_reg_10__12_ ( .D(add_fir[92]), .CK(clk), .Q(
        temp_add_fir[92]) );
  DFFQX1 temp_add_fir_reg_0__0_ ( .D(add_fir[240]), .CK(clk), .Q(
        temp_add_fir[237]) );
  DFFQX1 temp_add_fir_reg_10__10_ ( .D(add_fir[90]), .CK(clk), .Q(
        temp_add_fir[90]) );
  DFFQX1 temp_add_fir_reg_13__14_ ( .D(add_fir[46]), .CK(clk), .Q(
        temp_add_fir[46]) );
  DFFQX1 temp_add_fir_reg_9__11_ ( .D(add_fir[107]), .CK(clk), .Q(
        temp_add_fir[107]) );
  DFFQX2 temp_add_fir_reg_12__7_ ( .D(add_fir[55]), .CK(clk), .Q(
        temp_add_fir[55]) );
  DFFQX2 temp_add_fir_reg_12__8_ ( .D(add_fir[56]), .CK(clk), .Q(
        temp_add_fir[56]) );
  DFFQX2 temp_add_fir_reg_12__9_ ( .D(add_fir[57]), .CK(clk), .Q(
        temp_add_fir[57]) );
  DFFQX2 temp_add_fir_reg_15__13_ ( .D(add_fir[13]), .CK(clk), .Q(
        temp_add_fir[13]) );
  DFFQX2 temp_add_fir_reg_15__14_ ( .D(add_fir[14]), .CK(clk), .Q(
        temp_add_fir[14]) );
  DFFQX1 temp_mul_add_fir_reg_6__5_ ( .D(mul_add_fir[272]), .CK(clk), .Q(
        temp_mul_add_fir[293]) );
  DFFQX1 temp_mul_add_fir_reg_8__5_ ( .D(mul_add_fir[221]), .CK(clk), .Q(
        temp_mul_add_fir[229]) );
  DFFQX1 temp_mul_add_fir_reg_10__5_ ( .D(mul_add_fir[158]), .CK(clk), .Q(
        temp_mul_add_fir[165]) );
  DFFQX1 temp_mul_add_fir_reg_12__6_ ( .D(mul_add_fir[98]), .CK(clk), .Q(
        temp_mul_add_fir[102]) );
  DFFQX1 temp_mul_add_fir_reg_12__5_ ( .D(mul_add_fir[97]), .CK(clk), .Q(
        temp_mul_add_fir[101]) );
  DFFQX1 temp_add_fir_reg_13__9_ ( .D(add_fir[41]), .CK(clk), .Q(
        temp_add_fir[41]) );
  DFFQX1 temp_add_fir_reg_11__1_ ( .D(add_fir[65]), .CK(clk), .Q(
        temp_add_fir[65]) );
  DFFQX1 temp_add_fir_reg_3__1_ ( .D(add_fir[193]), .CK(clk), .Q(
        temp_add_fir[190]) );
  DFFQX1 temp_add_fir_reg_13__8_ ( .D(add_fir[40]), .CK(clk), .Q(
        temp_add_fir[40]) );
  DFFQX1 temp_mul_add_fir_reg_11__5_ ( .D(mul_add_fir[127]), .CK(clk), .Q(
        temp_mul_add_fir[133]) );
  DFFQX1 temp_add_fir_reg_2__1_ ( .D(add_fir[209]), .CK(clk), .Q(
        temp_add_fir[206]) );
  DFFQX1 temp_add_fir_reg_8__5_ ( .D(add_fir[117]), .CK(clk), .Q(
        temp_add_fir[117]) );
  DFFQX1 temp_add_fir_reg_9__4_ ( .D(add_fir[100]), .CK(clk), .Q(
        temp_add_fir[100]) );
  DFFQX1 temp_add_fir_reg_1__2_ ( .D(add_fir[226]), .CK(clk), .Q(
        temp_add_fir[223]) );
  DFFQX1 temp_add_fir_reg_11__3_ ( .D(add_fir[67]), .CK(clk), .Q(
        temp_add_fir[67]) );
  DFFQX1 temp_add_fir_reg_8__6_ ( .D(add_fir[118]), .CK(clk), .Q(
        temp_add_fir[118]) );
  DFFQX1 temp_add_fir_reg_8__7_ ( .D(add_fir[119]), .CK(clk), .Q(
        temp_add_fir[119]) );
  DFFQX1 temp_add_fir_reg_9__7_ ( .D(add_fir[103]), .CK(clk), .Q(
        temp_add_fir[103]) );
  DFFQX1 temp_add_fir_reg_9__6_ ( .D(add_fir[102]), .CK(clk), .Q(
        temp_add_fir[102]) );
  DFFQX1 temp_add_fir_reg_3__2_ ( .D(add_fir[194]), .CK(clk), .Q(
        temp_add_fir[191]) );
  DFFQX1 temp_add_fir_reg_2__2_ ( .D(add_fir[210]), .CK(clk), .Q(
        temp_add_fir[207]) );
  DFFQX1 temp_add_fir_reg_3__0_ ( .D(add_fir[192]), .CK(clk), .Q(
        temp_add_fir[189]) );
  DFFQX1 temp_add_fir_reg_11__2_ ( .D(add_fir[66]), .CK(clk), .Q(
        temp_add_fir[66]) );
  DFFQX1 temp_add_fir_reg_1__1_ ( .D(add_fir[225]), .CK(clk), .Q(
        temp_add_fir[222]) );
  DFFQX1 temp_add_fir_reg_10__6_ ( .D(add_fir[86]), .CK(clk), .Q(
        temp_add_fir[86]) );
  DFFQX1 temp_add_fir_reg_10__4_ ( .D(add_fir[84]), .CK(clk), .Q(
        temp_add_fir[84]) );
  DFFQX1 temp_add_fir_reg_2__3_ ( .D(add_fir[211]), .CK(clk), .Q(
        temp_add_fir[208]) );
  DFFQX1 temp_add_fir_reg_1__0_ ( .D(add_fir[224]), .CK(clk), .Q(
        temp_add_fir[221]) );
  DFFQX1 temp_add_fir_reg_10__5_ ( .D(add_fir[85]), .CK(clk), .Q(
        temp_add_fir[85]) );
  DFFQX1 temp_add_fir_reg_13__7_ ( .D(add_fir[39]), .CK(clk), .Q(
        temp_add_fir[39]) );
  DFFQX1 temp_add_fir_reg_8__4_ ( .D(add_fir[116]), .CK(clk), .Q(
        temp_add_fir[116]) );
  DFFQX1 temp_add_fir_reg_10__8_ ( .D(add_fir[88]), .CK(clk), .Q(
        temp_add_fir[88]) );
  DFFQX1 temp_add_fir_reg_9__5_ ( .D(add_fir[101]), .CK(clk), .Q(
        temp_add_fir[101]) );
  DFFQX1 temp_add_fir_reg_4__2_ ( .D(add_fir[178]), .CK(clk), .Q(
        temp_add_fir[175]) );
  DFFQX1 temp_add_fir_reg_4__3_ ( .D(add_fir[179]), .CK(clk), .Q(
        temp_add_fir[176]) );
  DFFQX1 temp_add_fir_reg_10__7_ ( .D(add_fir[87]), .CK(clk), .Q(
        temp_add_fir[87]) );
  DFFQX1 temp_add_fir_reg_4__0_ ( .D(add_fir[176]), .CK(clk), .Q(
        temp_add_fir[173]) );
  DFFQX1 temp_add_fir_reg_14__8_ ( .D(add_fir[24]), .CK(clk), .Q(
        temp_add_fir[24]) );
  DFFQX1 temp_add_fir_reg_12__0_ ( .D(add_fir[48]), .CK(clk), .Q(
        temp_add_fir[48]) );
  DFFQX1 temp_add_fir_reg_4__4_ ( .D(add_fir[180]), .CK(clk), .Q(
        temp_add_fir[177]) );
  DFFQX1 temp_add_fir_reg_4__1_ ( .D(add_fir[177]), .CK(clk), .Q(
        temp_add_fir[174]) );
  DFFQX1 temp_add_fir_reg_12__2_ ( .D(add_fir[50]), .CK(clk), .Q(
        temp_add_fir[50]) );
  DFFQX1 temp_add_fir_reg_14__6_ ( .D(add_fir[22]), .CK(clk), .Q(
        temp_add_fir[22]) );
  DFFQX1 temp_add_fir_reg_14__10_ ( .D(add_fir[26]), .CK(clk), .Q(
        temp_add_fir[26]) );
  DFFQX1 temp_add_fir_reg_12__1_ ( .D(add_fir[49]), .CK(clk), .Q(
        temp_add_fir[49]) );
  DFFQX1 temp_add_fir_reg_2__0_ ( .D(add_fir[208]), .CK(clk), .Q(
        temp_add_fir[205]) );
  DFFQX1 temp_add_fir_reg_12__3_ ( .D(add_fir[51]), .CK(clk), .Q(
        temp_add_fir[51]) );
  DFFQX2 temp_add_fir_reg_12__4_ ( .D(add_fir[52]), .CK(clk), .Q(
        temp_add_fir[52]) );
  DFFQX2 temp_add_fir_reg_11__0_ ( .D(add_fir[64]), .CK(clk), .Q(
        temp_add_fir[64]) );
  DFFQX2 temp_add_fir_reg_12__5_ ( .D(add_fir[53]), .CK(clk), .Q(
        temp_add_fir[53]) );
  DFFQX2 temp_add_fir_reg_12__6_ ( .D(add_fir[54]), .CK(clk), .Q(
        temp_add_fir[54]) );
  DFFQX2 temp_add_fir_reg_15__11_ ( .D(add_fir[11]), .CK(clk), .Q(
        temp_add_fir[11]) );
  DFFQX2 temp_add_fir_reg_15__9_ ( .D(add_fir[9]), .CK(clk), .Q(
        temp_add_fir[9]) );
  DFFQX2 temp_add_fir_reg_15__12_ ( .D(add_fir[12]), .CK(clk), .Q(
        temp_add_fir[12]) );
  DFFQX2 temp_add_fir_reg_15__10_ ( .D(add_fir[10]), .CK(clk), .Q(
        temp_add_fir[10]) );
  DFFQX1 temp_mul_add_fir_reg_0__4_ ( .D(mul_add_fir[460]), .CK(clk), .Q(
        temp_mul_add_fir[484]) );
  DFFQX1 temp_mul_add_fir_reg_0__3_ ( .D(mul_add_fir[459]), .CK(clk), .Q(
        temp_mul_add_fir[483]) );
  DFFQX1 temp_mul_add_fir_reg_0__2_ ( .D(mul_add_fir[458]), .CK(clk), .Q(
        temp_mul_add_fir[482]) );
  DFFQX1 temp_mul_add_fir_reg_2__4_ ( .D(mul_add_fir[398]), .CK(clk), .Q(
        temp_mul_add_fir[420]) );
  DFFQX1 temp_mul_add_fir_reg_2__3_ ( .D(mul_add_fir[397]), .CK(clk), .Q(
        temp_mul_add_fir[419]) );
  DFFQX1 temp_mul_add_fir_reg_2__2_ ( .D(mul_add_fir[396]), .CK(clk), .Q(
        temp_mul_add_fir[418]) );
  DFFQX1 temp_mul_add_fir_reg_4__4_ ( .D(mul_add_fir[334]), .CK(clk), .Q(
        temp_mul_add_fir[356]) );
  DFFQX1 temp_mul_add_fir_reg_4__2_ ( .D(mul_add_fir[332]), .CK(clk), .Q(
        temp_mul_add_fir[354]) );
  DFFQX1 temp_mul_add_fir_reg_6__4_ ( .D(mul_add_fir[271]), .CK(clk), .Q(
        temp_mul_add_fir[292]) );
  DFFQX1 temp_mul_add_fir_reg_6__3_ ( .D(mul_add_fir[270]), .CK(clk), .Q(
        temp_mul_add_fir[291]) );
  DFFQX1 temp_mul_add_fir_reg_6__2_ ( .D(mul_add_fir[269]), .CK(clk), .Q(
        temp_mul_add_fir[290]) );
  DFFQX1 temp_mul_add_fir_reg_8__4_ ( .D(mul_add_fir[220]), .CK(clk), .Q(
        temp_mul_add_fir[228]) );
  DFFQX1 temp_mul_add_fir_reg_8__3_ ( .D(mul_add_fir[219]), .CK(clk), .Q(
        temp_mul_add_fir[227]) );
  DFFQX1 temp_mul_add_fir_reg_8__2_ ( .D(mul_add_fir[218]), .CK(clk), .Q(
        temp_mul_add_fir[226]) );
  DFFQX1 temp_mul_add_fir_reg_10__4_ ( .D(mul_add_fir[157]), .CK(clk), .Q(
        temp_mul_add_fir[164]) );
  DFFQX1 temp_mul_add_fir_reg_10__3_ ( .D(mul_add_fir[156]), .CK(clk), .Q(
        temp_mul_add_fir[163]) );
  DFFQX1 temp_mul_add_fir_reg_10__2_ ( .D(mul_add_fir[155]), .CK(clk), .Q(
        temp_mul_add_fir[162]) );
  DFFQX1 temp_mul_add_fir_reg_12__4_ ( .D(mul_add_fir[96]), .CK(clk), .Q(
        temp_mul_add_fir[100]) );
  DFFQX1 temp_mul_add_fir_reg_12__3_ ( .D(mul_add_fir[95]), .CK(clk), .Q(
        temp_mul_add_fir[99]) );
  DFFQX1 temp_mul_add_fir_reg_12__2_ ( .D(mul_add_fir[94]), .CK(clk), .Q(
        temp_mul_add_fir[98]) );
  DFFQX1 temp_mul_add_fir_reg_14__4_ ( .D(mul_add_fir[35]), .CK(clk), .Q(
        temp_mul_add_fir[36]) );
  DFFQX1 temp_mul_add_fir_reg_14__3_ ( .D(mul_add_fir[34]), .CK(clk), .Q(
        temp_mul_add_fir[35]) );
  DFFQX1 temp_mul_add_fir_reg_14__2_ ( .D(mul_add_fir[33]), .CK(clk), .Q(
        temp_mul_add_fir[34]) );
  DFFQX1 temp_add_fir_reg_13__6_ ( .D(add_fir[38]), .CK(clk), .Q(
        temp_add_fir[38]) );
  DFFQX1 temp_add_fir_reg_13__5_ ( .D(add_fir[37]), .CK(clk), .Q(
        temp_add_fir[37]) );
  DFFQX1 temp_add_fir_reg_13__3_ ( .D(add_fir[35]), .CK(clk), .Q(
        temp_add_fir[35]) );
  DFFQX1 temp_add_fir_reg_13__1_ ( .D(add_fir[33]), .CK(clk), .Q(
        temp_add_fir[33]) );
  DFFQX1 temp_mul_add_fir_reg_1__4_ ( .D(mul_add_fir[429]), .CK(clk), .Q(
        temp_mul_add_fir[452]) );
  DFFQX1 temp_mul_add_fir_reg_1__3_ ( .D(mul_add_fir[428]), .CK(clk), .Q(
        temp_mul_add_fir[451]) );
  DFFQX1 temp_mul_add_fir_reg_1__2_ ( .D(mul_add_fir[427]), .CK(clk), .Q(
        temp_mul_add_fir[450]) );
  DFFQX1 temp_mul_add_fir_reg_3__4_ ( .D(mul_add_fir[366]), .CK(clk), .Q(
        temp_mul_add_fir[388]) );
  DFFQX1 temp_mul_add_fir_reg_3__3_ ( .D(mul_add_fir[365]), .CK(clk), .Q(
        temp_mul_add_fir[387]) );
  DFFQX1 temp_mul_add_fir_reg_3__2_ ( .D(mul_add_fir[364]), .CK(clk), .Q(
        temp_mul_add_fir[386]) );
  DFFQX1 temp_mul_add_fir_reg_5__4_ ( .D(mul_add_fir[302]), .CK(clk), .Q(
        temp_mul_add_fir[324]) );
  DFFQX1 temp_mul_add_fir_reg_5__2_ ( .D(mul_add_fir[300]), .CK(clk), .Q(
        temp_mul_add_fir[322]) );
  DFFQX1 temp_mul_add_fir_reg_7__4_ ( .D(mul_add_fir[250]), .CK(clk), .Q(
        temp_mul_add_fir[260]) );
  DFFQX1 temp_mul_add_fir_reg_7__3_ ( .D(mul_add_fir[249]), .CK(clk), .Q(
        temp_mul_add_fir[259]) );
  DFFQX1 temp_mul_add_fir_reg_7__2_ ( .D(mul_add_fir[248]), .CK(clk), .Q(
        temp_mul_add_fir[258]) );
  DFFQX1 temp_mul_add_fir_reg_9__4_ ( .D(mul_add_fir[188]), .CK(clk), .Q(
        temp_mul_add_fir[196]) );
  DFFQX1 temp_mul_add_fir_reg_9__3_ ( .D(mul_add_fir[187]), .CK(clk), .Q(
        temp_mul_add_fir[195]) );
  DFFQX1 temp_mul_add_fir_reg_9__2_ ( .D(mul_add_fir[186]), .CK(clk), .Q(
        temp_mul_add_fir[194]) );
  DFFQX1 temp_mul_add_fir_reg_11__4_ ( .D(mul_add_fir[126]), .CK(clk), .Q(
        temp_mul_add_fir[132]) );
  DFFQX1 temp_mul_add_fir_reg_11__3_ ( .D(mul_add_fir[125]), .CK(clk), .Q(
        temp_mul_add_fir[131]) );
  DFFQX1 temp_mul_add_fir_reg_11__2_ ( .D(mul_add_fir[124]), .CK(clk), .Q(
        temp_mul_add_fir[130]) );
  DFFQX1 temp_mul_add_fir_reg_13__4_ ( .D(mul_add_fir[65]), .CK(clk), .Q(
        temp_mul_add_fir[68]) );
  DFFQX1 temp_mul_add_fir_reg_13__3_ ( .D(mul_add_fir[64]), .CK(clk), .Q(
        temp_mul_add_fir[67]) );
  DFFQX1 temp_mul_add_fir_reg_13__2_ ( .D(mul_add_fir[63]), .CK(clk), .Q(
        temp_mul_add_fir[66]) );
  DFFQX1 temp_mul_add_fir_reg_15__4_ ( .D(mul_add_fir[4]), .CK(clk), .Q(
        temp_mul_add_fir[4]) );
  DFFQX1 temp_mul_add_fir_reg_15__3_ ( .D(mul_add_fir[3]), .CK(clk), .Q(
        temp_mul_add_fir[3]) );
  DFFQX1 temp_mul_add_fir_reg_15__2_ ( .D(mul_add_fir[2]), .CK(clk), .Q(
        temp_mul_add_fir[2]) );
  DFFQX1 temp_add_fir_reg_10__1_ ( .D(add_fir[81]), .CK(clk), .Q(
        temp_add_fir[81]) );
  DFFQX1 temp_add_fir_reg_8__3_ ( .D(add_fir[115]), .CK(clk), .Q(
        temp_add_fir[115]) );
  DFFQX1 temp_add_fir_reg_9__3_ ( .D(add_fir[99]), .CK(clk), .Q(
        temp_add_fir[99]) );
  DFFQX1 temp_add_fir_reg_8__1_ ( .D(add_fir[113]), .CK(clk), .Q(
        temp_add_fir[113]) );
  DFFQX1 temp_add_fir_reg_9__1_ ( .D(add_fir[97]), .CK(clk), .Q(
        temp_add_fir[97]) );
  DFFQX1 temp_add_fir_reg_13__4_ ( .D(add_fir[36]), .CK(clk), .Q(
        temp_add_fir[36]) );
  DFFQX1 temp_add_fir_reg_13__2_ ( .D(add_fir[34]), .CK(clk), .Q(
        temp_add_fir[34]) );
  DFFQX1 temp_add_fir_reg_10__2_ ( .D(add_fir[82]), .CK(clk), .Q(
        temp_add_fir[82]) );
  DFFQX1 temp_add_fir_reg_13__0_ ( .D(add_fir[32]), .CK(clk), .Q(
        temp_add_fir[32]) );
  DFFQX1 temp_add_fir_reg_8__2_ ( .D(add_fir[114]), .CK(clk), .Q(
        temp_add_fir[114]) );
  DFFQX1 temp_add_fir_reg_9__2_ ( .D(add_fir[98]), .CK(clk), .Q(
        temp_add_fir[98]) );
  DFFQX1 temp_add_fir_reg_14__2_ ( .D(add_fir[18]), .CK(clk), .Q(
        temp_add_fir[18]) );
  DFFQX1 temp_add_fir_reg_14__4_ ( .D(add_fir[20]), .CK(clk), .Q(
        temp_add_fir[20]) );
  DFFQX1 temp_add_fir_reg_14__3_ ( .D(add_fir[19]), .CK(clk), .Q(
        temp_add_fir[19]) );
  DFFQX1 temp_add_fir_reg_14__1_ ( .D(add_fir[17]), .CK(clk), .Q(
        temp_add_fir[17]) );
  DFFQX1 temp_add_fir_reg_14__7_ ( .D(add_fir[23]), .CK(clk), .Q(
        temp_add_fir[23]) );
  DFFQX1 temp_add_fir_reg_14__5_ ( .D(add_fir[21]), .CK(clk), .Q(
        temp_add_fir[21]) );
  DFFQX1 temp_add_fir_reg_10__3_ ( .D(add_fir[83]), .CK(clk), .Q(
        temp_add_fir[83]) );
  DFFQX1 temp_add_fir_reg_8__0_ ( .D(add_fir[112]), .CK(clk), .Q(
        temp_add_fir[112]) );
  DFFQX1 temp_add_fir_reg_9__0_ ( .D(add_fir[96]), .CK(clk), .Q(
        temp_add_fir[96]) );
  DFFQX1 temp_add_fir_reg_10__0_ ( .D(add_fir[80]), .CK(clk), .Q(
        temp_add_fir[80]) );
  DFFQX2 temp_add_fir_reg_15__4_ ( .D(add_fir[4]), .CK(clk), .Q(
        temp_add_fir[4]) );
  DFFQX2 temp_add_fir_reg_15__0_ ( .D(add_fir[0]), .CK(clk), .Q(
        temp_add_fir[0]) );
  DFFQX2 temp_add_fir_reg_15__3_ ( .D(add_fir[3]), .CK(clk), .Q(
        temp_add_fir[3]) );
  DFFQX2 temp_add_fir_reg_15__7_ ( .D(add_fir[7]), .CK(clk), .Q(
        temp_add_fir[7]) );
  DFFQX2 temp_add_fir_reg_14__0_ ( .D(add_fir[16]), .CK(clk), .Q(
        temp_add_fir[16]) );
  DFFQX2 temp_add_fir_reg_15__1_ ( .D(add_fir[1]), .CK(clk), .Q(
        temp_add_fir[1]) );
  DFFQX2 temp_add_fir_reg_15__6_ ( .D(add_fir[6]), .CK(clk), .Q(
        temp_add_fir[6]) );
  DFFQX2 temp_add_fir_reg_15__5_ ( .D(add_fir[5]), .CK(clk), .Q(
        temp_add_fir[5]) );
  DFFQX2 temp_add_fir_reg_15__8_ ( .D(add_fir[8]), .CK(clk), .Q(
        temp_add_fir[8]) );
  DFFQX1 temp_mul_add_fir_reg_0__1_ ( .D(mul_add_fir[457]), .CK(clk), .Q(
        temp_mul_add_fir[481]) );
  DFFQX1 temp_mul_add_fir_reg_2__1_ ( .D(mul_add_fir[395]), .CK(clk), .Q(
        temp_mul_add_fir[417]) );
  DFFQX1 temp_mul_add_fir_reg_4__1_ ( .D(mul_add_fir[331]), .CK(clk), .Q(
        temp_mul_add_fir[353]) );
  DFFQX1 temp_mul_add_fir_reg_6__1_ ( .D(mul_add_fir[268]), .CK(clk), .Q(
        temp_mul_add_fir[289]) );
  DFFQX1 temp_mul_add_fir_reg_8__1_ ( .D(mul_add_fir[217]), .CK(clk), .Q(
        temp_mul_add_fir[225]) );
  DFFQX1 temp_mul_add_fir_reg_10__1_ ( .D(mul_add_fir[154]), .CK(clk), .Q(
        temp_mul_add_fir[161]) );
  DFFQX1 temp_mul_add_fir_reg_12__1_ ( .D(mul_add_fir[93]), .CK(clk), .Q(
        temp_mul_add_fir[97]) );
  DFFQX1 temp_mul_add_fir_reg_14__1_ ( .D(mul_add_fir[32]), .CK(clk), .Q(
        temp_mul_add_fir[33]) );
  DFFQX1 temp_mul_add_fir_reg_1__1_ ( .D(mul_add_fir[426]), .CK(clk), .Q(
        temp_mul_add_fir[449]) );
  DFFQX1 temp_mul_add_fir_reg_3__1_ ( .D(mul_add_fir[363]), .CK(clk), .Q(
        temp_mul_add_fir[385]) );
  DFFQX1 temp_mul_add_fir_reg_5__1_ ( .D(mul_add_fir[299]), .CK(clk), .Q(
        temp_mul_add_fir[321]) );
  DFFQX1 temp_mul_add_fir_reg_9__1_ ( .D(mul_add_fir[185]), .CK(clk), .Q(
        temp_mul_add_fir[193]) );
  DFFQX1 temp_mul_add_fir_reg_15__1_ ( .D(mul_add_fir[1]), .CK(clk), .Q(
        temp_mul_add_fir[1]) );
  ADDHXL add_55_U1_1_4 ( .A(cnt_data[4]), .B(add_55_carry[4]), .CO(
        add_55_carry[5]), .S(N16) );
  ADDHXL add_55_U1_1_3 ( .A(cnt_data[3]), .B(add_55_carry[3]), .CO(
        add_55_carry[4]), .S(N15) );
  ADDHXL add_55_U1_1_2 ( .A(cnt_data[2]), .B(add_55_carry[2]), .CO(
        add_55_carry[3]), .S(N14) );
  ADDHXL add_55_U1_1_1 ( .A(cnt_data[1]), .B(cnt_data[0]), .CO(add_55_carry[2]), .S(N13) );
  DFFRX1 cnt_data_reg_1_ ( .D(n1020), .CK(clk), .RN(n1030), .Q(cnt_data[1]), 
        .QN(n58) );
  DFFQX1 temp_add_fir_reg_14__9_ ( .D(add_fir[25]), .CK(clk), .Q(
        temp_add_fir[25]) );
  DFFQX1 temp_add_fir_reg_15__2_ ( .D(add_fir[2]), .CK(clk), .Q(
        temp_add_fir[2]) );
  DFFQX1 temp_mul_add_fir_reg_10__8_ ( .D(mul_add_fir[161]), .CK(clk), .Q(
        temp_mul_add_fir[168]) );
  DFFQX1 temp_mul_add_fir_reg_9__8_ ( .D(mul_add_fir[192]), .CK(clk), .Q(
        temp_mul_add_fir[200]) );
  DFFQX1 temp_mul_add_fir_reg_11__8_ ( .D(mul_add_fir[130]), .CK(clk), .Q(
        temp_mul_add_fir[136]) );
  DFFQX1 temp_mul_add_fir_reg_2__8_ ( .D(mul_add_fir[402]), .CK(clk), .Q(
        temp_mul_add_fir[424]) );
  DFFQX1 temp_mul_add_fir_reg_4__7_ ( .D(mul_add_fir[337]), .CK(clk), .Q(
        temp_mul_add_fir[359]) );
  DFFQX1 temp_mul_add_fir_reg_8__6_ ( .D(mul_add_fir[222]), .CK(clk), .Q(
        temp_mul_add_fir[230]) );
  DFFQX1 temp_mul_add_fir_reg_14__7_ ( .D(mul_add_fir[38]), .CK(clk), .Q(
        temp_mul_add_fir[39]) );
  DFFQX1 temp_mul_add_fir_reg_3__8_ ( .D(mul_add_fir[370]), .CK(clk), .Q(
        temp_mul_add_fir[392]) );
  DFFQX1 temp_mul_add_fir_reg_5__7_ ( .D(mul_add_fir[305]), .CK(clk), .Q(
        temp_mul_add_fir[327]) );
  DFFQX1 temp_mul_add_fir_reg_15__7_ ( .D(mul_add_fir[7]), .CK(clk), .Q(
        temp_mul_add_fir[7]) );
  DFFQX1 temp_mul_add_fir_reg_10__7_ ( .D(mul_add_fir[160]), .CK(clk), .Q(
        temp_mul_add_fir[167]) );
  DFFQX1 temp_mul_add_fir_reg_12__7_ ( .D(mul_add_fir[99]), .CK(clk), .Q(
        temp_mul_add_fir[103]) );
  DFFQX1 temp_mul_add_fir_reg_6__8_ ( .D(mul_add_fir[275]), .CK(clk), .Q(
        temp_mul_add_fir[296]) );
  DFFQX1 temp_mul_add_fir_reg_6__7_ ( .D(mul_add_fir[274]), .CK(clk), .Q(
        temp_mul_add_fir[295]) );
  DFFQX1 temp_mul_add_fir_reg_7__8_ ( .D(mul_add_fir[254]), .CK(clk), .Q(
        temp_mul_add_fir[264]) );
  DFFQX1 temp_mul_add_fir_reg_7__7_ ( .D(mul_add_fir[253]), .CK(clk), .Q(
        temp_mul_add_fir[263]) );
  DFFQX1 temp_mul_add_fir_reg_13__8_ ( .D(mul_add_fir[69]), .CK(clk), .Q(
        temp_mul_add_fir[72]) );
  DFFQX1 temp_mul_add_fir_reg_8__7_ ( .D(mul_add_fir[223]), .CK(clk), .Q(
        temp_mul_add_fir[231]) );
  DFFQX1 temp_mul_add_fir_reg_14__8_ ( .D(mul_add_fir[39]), .CK(clk), .Q(
        temp_mul_add_fir[40]) );
  DFFQX1 temp_mul_add_fir_reg_11__7_ ( .D(mul_add_fir[129]), .CK(clk), .Q(
        temp_mul_add_fir[135]) );
  DFFQX1 temp_mul_add_fir_reg_13__7_ ( .D(mul_add_fir[68]), .CK(clk), .Q(
        temp_mul_add_fir[71]) );
  DFFQX1 temp_mul_add_fir_reg_5__8_ ( .D(mul_add_fir[306]), .CK(clk), .Q(
        temp_mul_add_fir[328]) );
  DFFQX1 temp_mul_add_fir_reg_9__7_ ( .D(mul_add_fir[191]), .CK(clk), .Q(
        temp_mul_add_fir[199]) );
  DFFQX1 temp_mul_add_fir_reg_15__8_ ( .D(mul_add_fir[8]), .CK(clk), .Q(
        temp_mul_add_fir[8]) );
  DFFRX2 fir_d_reg_15_ ( .D(revise_o[15]), .CK(clk), .RN(n1030), .QN(n33) );
  DFFRX1 cnt_data_reg_3_ ( .D(n1000), .CK(clk), .RN(n1030), .Q(cnt_data[3]), 
        .QN(n940) );
  DFFRX1 cnt_data_reg_4_ ( .D(n990), .CK(clk), .RN(n1030), .Q(cnt_data[4]) );
  DFFRX1 cnt_data_reg_2_ ( .D(n1010), .CK(clk), .RN(n1030), .Q(cnt_data[2]) );
  DFFRX1 cnt_data_reg_5_ ( .D(n980), .CK(clk), .RN(n1030), .Q(cnt_data[5]) );
  DFFRX1 cnt_data_reg_0_ ( .D(n970), .CK(clk), .RN(n1030), .Q(cnt_data[0]), 
        .QN(N12) );
  DFFSRHQX1 fir_valid_state_reg ( .D(N54), .CK(clk), .SN(1'b1), .RN(n1030), 
        .Q(n149) );
  DFFQX1 temp_mul_add_fir_reg_10__6_ ( .D(mul_add_fir[159]), .CK(clk), .Q(
        temp_mul_add_fir[166]) );
  DFFQX1 temp_mul_add_fir_reg_14__6_ ( .D(mul_add_fir[37]), .CK(clk), .Q(
        temp_mul_add_fir[38]) );
  DFFQX1 temp_mul_add_fir_reg_0__6_ ( .D(mul_add_fir[462]), .CK(clk), .Q(
        temp_mul_add_fir[486]) );
  DFFQX1 temp_mul_add_fir_reg_4__6_ ( .D(mul_add_fir[336]), .CK(clk), .Q(
        temp_mul_add_fir[358]) );
  DFFQX1 temp_mul_add_fir_reg_0__7_ ( .D(mul_add_fir[463]), .CK(clk), .Q(
        temp_mul_add_fir[487]) );
  DFFQX1 temp_mul_add_fir_reg_2__6_ ( .D(mul_add_fir[400]), .CK(clk), .Q(
        temp_mul_add_fir[422]) );
  DFFQX1 temp_mul_add_fir_reg_2__7_ ( .D(mul_add_fir[401]), .CK(clk), .Q(
        temp_mul_add_fir[423]) );
  DFFQX1 temp_mul_add_fir_reg_11__6_ ( .D(mul_add_fir[128]), .CK(clk), .Q(
        temp_mul_add_fir[134]) );
  DFFQX1 temp_mul_add_fir_reg_13__6_ ( .D(mul_add_fir[67]), .CK(clk), .Q(
        temp_mul_add_fir[70]) );
  DFFQX1 temp_mul_add_fir_reg_1__6_ ( .D(mul_add_fir[431]), .CK(clk), .Q(
        temp_mul_add_fir[454]) );
  DFFQX1 temp_mul_add_fir_reg_9__6_ ( .D(mul_add_fir[190]), .CK(clk), .Q(
        temp_mul_add_fir[198]) );
  DFFQX1 temp_mul_add_fir_reg_3__6_ ( .D(mul_add_fir[368]), .CK(clk), .Q(
        temp_mul_add_fir[390]) );
  DFFQX1 temp_mul_add_fir_reg_1__7_ ( .D(mul_add_fir[432]), .CK(clk), .Q(
        temp_mul_add_fir[455]) );
  DFFQX1 temp_mul_add_fir_reg_3__7_ ( .D(mul_add_fir[369]), .CK(clk), .Q(
        temp_mul_add_fir[391]) );
  DFFQX1 temp_mul_add_fir_reg_14__5_ ( .D(mul_add_fir[36]), .CK(clk), .Q(
        temp_mul_add_fir[37]) );
  DFFQX1 temp_mul_add_fir_reg_4__5_ ( .D(mul_add_fir[335]), .CK(clk), .Q(
        temp_mul_add_fir[357]) );
  DFFQX1 temp_mul_add_fir_reg_0__5_ ( .D(mul_add_fir[461]), .CK(clk), .Q(
        temp_mul_add_fir[485]) );
  DFFQX1 temp_mul_add_fir_reg_2__5_ ( .D(mul_add_fir[399]), .CK(clk), .Q(
        temp_mul_add_fir[421]) );
  DFFQX1 temp_mul_add_fir_reg_6__6_ ( .D(mul_add_fir[273]), .CK(clk), .Q(
        temp_mul_add_fir[294]) );
  DFFQX1 temp_mul_add_fir_reg_7__5_ ( .D(mul_add_fir[251]), .CK(clk), .Q(
        temp_mul_add_fir[261]) );
  DFFQX1 temp_mul_add_fir_reg_13__5_ ( .D(mul_add_fir[66]), .CK(clk), .Q(
        temp_mul_add_fir[69]) );
  DFFQX1 temp_mul_add_fir_reg_15__5_ ( .D(mul_add_fir[5]), .CK(clk), .Q(
        temp_mul_add_fir[5]) );
  DFFQX1 temp_mul_add_fir_reg_9__5_ ( .D(mul_add_fir[189]), .CK(clk), .Q(
        temp_mul_add_fir[197]) );
  DFFQX1 temp_mul_add_fir_reg_5__5_ ( .D(mul_add_fir[303]), .CK(clk), .Q(
        temp_mul_add_fir[325]) );
  DFFQX1 temp_mul_add_fir_reg_1__5_ ( .D(mul_add_fir[430]), .CK(clk), .Q(
        temp_mul_add_fir[453]) );
  DFFQX1 temp_mul_add_fir_reg_3__5_ ( .D(mul_add_fir[367]), .CK(clk), .Q(
        temp_mul_add_fir[389]) );
  DFFQX1 temp_mul_add_fir_reg_7__6_ ( .D(mul_add_fir[252]), .CK(clk), .Q(
        temp_mul_add_fir[262]) );
  DFFQX1 temp_mul_add_fir_reg_15__6_ ( .D(mul_add_fir[6]), .CK(clk), .Q(
        temp_mul_add_fir[6]) );
  DFFQX1 temp_mul_add_fir_reg_5__6_ ( .D(mul_add_fir[304]), .CK(clk), .Q(
        temp_mul_add_fir[326]) );
  DFFQX1 temp_mul_add_fir_reg_8__0_ ( .D(mul_add_fir[216]), .CK(clk), .Q(
        temp_mul_add_fir[224]) );
  DFFQX1 temp_mul_add_fir_reg_4__0_ ( .D(mul_add_fir[330]), .CK(clk), .Q(
        temp_mul_add_fir[352]) );
  DFFQX1 temp_mul_add_fir_reg_15__0_ ( .D(mul_add_fir[0]), .CK(clk), .Q(
        temp_mul_add_fir[0]) );
  DFFQX1 temp_mul_add_fir_reg_2__0_ ( .D(mul_add_fir[394]), .CK(clk), .Q(
        temp_mul_add_fir[416]) );
  DFFQX1 temp_mul_add_fir_reg_3__0_ ( .D(mul_add_fir[362]), .CK(clk), .Q(
        temp_mul_add_fir[384]) );
  DFFQX2 temp_mul_add_fir_reg_5__3_ ( .D(mul_add_fir[301]), .CK(clk), .Q(
        temp_mul_add_fir[323]) );
  DFFQX2 temp_mul_add_fir_reg_4__3_ ( .D(mul_add_fir[333]), .CK(clk), .Q(
        temp_mul_add_fir[355]) );
  INVX6 U4 ( .A(n540), .Y(n960) );
  BUFX12 U5 ( .A(comb_fir_o[31]), .Y(n540) );
  INVX16 U22 ( .A(n18), .Y(fir_d[0]) );
  INVX16 U23 ( .A(n19), .Y(fir_d[1]) );
  INVX16 U24 ( .A(n2010), .Y(fir_d[2]) );
  INVX16 U25 ( .A(n2110), .Y(fir_d[3]) );
  INVX16 U26 ( .A(n2410), .Y(fir_d[4]) );
  INVX16 U27 ( .A(n25), .Y(fir_d[5]) );
  NOR3XL U28 ( .A(cnt_data[2]), .B(cnt_data[4]), .C(cnt_data[3]), .Y(n61) );
  XNOR2XL U29 ( .A(cnt_data[4]), .B(n920), .Y(N23) );
  NOR2XL U30 ( .A(cnt_data[4]), .B(n920), .Y(n930) );
  NAND4XL U31 ( .A(cnt_data[1]), .B(cnt_data[0]), .C(cnt_data[5]), .D(n61), 
        .Y(n60) );
  XOR2XL U32 ( .A(add_55_carry[5]), .B(cnt_data[5]), .Y(N17) );
  XOR2XL U33 ( .A(cnt_data[5]), .B(n930), .Y(N24) );
  AOI22XL U34 ( .A0(cnt_data[5]), .A1(cnt_data[4]), .B0(n950), .B1(cnt_data[5]), .Y(N7) );
  OR2XL U35 ( .A(cnt_data[5]), .B(cnt_data[4]), .Y(n72) );
  INVX16 U36 ( .A(n2310), .Y(fir_d[6]) );
  INVX16 U37 ( .A(n2210), .Y(fir_d[7]) );
  INVX16 U38 ( .A(n26), .Y(fir_d[8]) );
  INVX16 U39 ( .A(n27), .Y(fir_d[9]) );
  INVX16 U40 ( .A(n28), .Y(fir_d[10]) );
  INVX16 U41 ( .A(n29), .Y(fir_d[11]) );
  INVX16 U42 ( .A(n30), .Y(fir_d[12]) );
  INVX16 U43 ( .A(n31), .Y(fir_d[13]) );
  INVX16 U44 ( .A(n32), .Y(fir_d[14]) );
  INVX16 U45 ( .A(n33), .Y(fir_d[15]) );
  CLKINVX1 U46 ( .A(n149), .Y(n50) );
  INVX16 U47 ( .A(n50), .Y(fir_valid) );
  AO22X1 U49 ( .A0(comb_fir_o[17]), .A1(n960), .B0(N506), .B1(n540), .Y(
        revise_o[1]) );
  AO22XL U50 ( .A0(comb_fir_o[19]), .A1(n960), .B0(N508), .B1(n540), .Y(
        revise_o[3]) );
  AO22XL U51 ( .A0(comb_fir_o[20]), .A1(n960), .B0(N509), .B1(n540), .Y(
        revise_o[4]) );
  AO22XL U52 ( .A0(comb_fir_o[21]), .A1(n960), .B0(N510), .B1(n540), .Y(
        revise_o[5]) );
  AO22XL U53 ( .A0(comb_fir_o[18]), .A1(n960), .B0(N507), .B1(n540), .Y(
        revise_o[2]) );
  INVX4 U54 ( .A(n540), .Y(n53) );
  AO22XL U55 ( .A0(comb_fir_o[16]), .A1(n960), .B0(N505), .B1(n540), .Y(
        revise_o[0]) );
  CLKBUFX3 U56 ( .A(temp_add_fir[63]), .Y(n570) );
  AO22X1 U57 ( .A0(comb_fir_o[25]), .A1(n960), .B0(n540), .B1(N514), .Y(
        revise_o[9]) );
  AO22X1 U58 ( .A0(comb_fir_o[22]), .A1(n53), .B0(N511), .B1(n540), .Y(
        revise_o[6]) );
  AO22X1 U59 ( .A0(comb_fir_o[23]), .A1(n53), .B0(N512), .B1(n540), .Y(
        revise_o[7]) );
  AO22X1 U60 ( .A0(comb_fir_o[24]), .A1(n53), .B0(N513), .B1(n540), .Y(
        revise_o[8]) );
  AO22X1 U61 ( .A0(comb_fir_o[26]), .A1(n53), .B0(N515), .B1(n540), .Y(
        revise_o[10]) );
  AO22X1 U62 ( .A0(comb_fir_o[27]), .A1(n53), .B0(N516), .B1(n540), .Y(
        revise_o[11]) );
  AO22X1 U63 ( .A0(comb_fir_o[28]), .A1(n53), .B0(N517), .B1(n540), .Y(
        revise_o[12]) );
  AO22X1 U64 ( .A0(comb_fir_o[29]), .A1(n53), .B0(N518), .B1(n540), .Y(
        revise_o[13]) );
  AO22X1 U65 ( .A0(comb_fir_o[30]), .A1(n53), .B0(N519), .B1(n540), .Y(
        revise_o[14]) );
  AND2X2 U66 ( .A(N520), .B(n540), .Y(revise_o[15]) );
  NOR2BX1 U67 ( .AN(n56), .B(n64), .Y(n66) );
  CLKBUFX3 U68 ( .A(mul_add_fir[267]), .Y(n55) );
  CLKINVX1 U69 ( .A(mult_120_n14), .Y(mul_add_fir[267]) );
  AOI2BB1X2 U70 ( .A0N(cnt_data[1]), .A1N(n62), .B0(n56), .Y(n65) );
  CLKINVX1 U71 ( .A(temp_add_fir[139]), .Y(n880) );
  CLKINVX1 U72 ( .A(n69), .Y(n1010) );
  AOI222XL U73 ( .A0(N14), .A1(n64), .B0(N21), .B1(n65), .C0(cnt_data[2]), 
        .C1(n66), .Y(n69) );
  CLKINVX1 U74 ( .A(n67), .Y(n990) );
  AOI222XL U75 ( .A0(N16), .A1(n64), .B0(N23), .B1(n65), .C0(cnt_data[4]), 
        .C1(n66), .Y(n67) );
  CLKINVX1 U76 ( .A(temp_add_fir[137]), .Y(n860) );
  CLKINVX1 U77 ( .A(temp_add_fir[140]), .Y(n890) );
  CLKINVX1 U78 ( .A(temp_add_fir[138]), .Y(n870) );
  CLKINVX1 U79 ( .A(mul_add_fir[249]), .Y(n750) );
  CLKINVX1 U80 ( .A(mul_add_fir[250]), .Y(n760) );
  CLKINVX1 U81 ( .A(temp_add_fir[129]), .Y(n780) );
  CLKINVX1 U82 ( .A(temp_add_fir[130]), .Y(n790) );
  CLKINVX1 U83 ( .A(temp_add_fir[131]), .Y(n800) );
  CLKINVX1 U84 ( .A(temp_add_fir[132]), .Y(n810) );
  CLKINVX1 U85 ( .A(temp_add_fir[133]), .Y(n820) );
  CLKINVX1 U86 ( .A(temp_add_fir[134]), .Y(n830) );
  CLKINVX1 U87 ( .A(temp_add_fir[135]), .Y(n840) );
  CLKINVX1 U88 ( .A(temp_add_fir[136]), .Y(n850) );
  AND2X2 U89 ( .A(N7), .B(n56), .Y(n64) );
  CLKBUFX3 U90 ( .A(data_valid), .Y(n56) );
  CLKINVX1 U91 ( .A(n71), .Y(n970) );
  AOI222XL U92 ( .A0(N12), .A1(n64), .B0(N12), .B1(n65), .C0(n66), .C1(
        cnt_data[0]), .Y(n71) );
  CLKINVX1 U93 ( .A(n68), .Y(n1000) );
  AOI222XL U94 ( .A0(N15), .A1(n64), .B0(N22), .B1(n65), .C0(cnt_data[3]), 
        .C1(n66), .Y(n68) );
  CLKINVX1 U95 ( .A(n63), .Y(n980) );
  AOI222XL U96 ( .A0(N17), .A1(n64), .B0(N24), .B1(n65), .C0(n66), .C1(
        cnt_data[5]), .Y(n63) );
  CLKINVX1 U97 ( .A(n701), .Y(n1020) );
  AOI222XL U98 ( .A0(N13), .A1(n64), .B0(N20), .B1(n65), .C0(n66), .C1(
        cnt_data[1]), .Y(n701) );
  CLKINVX1 U99 ( .A(temp_add_fir[128]), .Y(n770) );
  CLKBUFX3 U100 ( .A(temp_add_fir[156]), .Y(n730) );
  CLKBUFX3 U101 ( .A(temp_add_fir[172]), .Y(n740) );
  OR2X1 U102 ( .A(cnt_data[1]), .B(cnt_data[0]), .Y(n900) );
  NAND2X1 U103 ( .A(n59), .B(n60), .Y(N54) );
  OAI21XL U104 ( .A0(n58), .A1(n62), .B0(fir_valid), .Y(n59) );
  OR4X1 U105 ( .A(cnt_data[0]), .B(cnt_data[2]), .C(n72), .D(cnt_data[3]), .Y(
        n62) );
  NAND2X1 U120 ( .A(mul_add_fir[248]), .B(n770), .Y(mult_120_n29) );
  XOR2X1 U121 ( .A(temp_add_fir[128]), .B(mul_add_fir[248]), .Y(
        mul_add_fir[251]) );
  OAI2BB1X1 U122 ( .A0N(cnt_data[0]), .A1N(cnt_data[1]), .B0(n900), .Y(N20) );
  NOR2X1 U123 ( .A(n900), .B(cnt_data[2]), .Y(n910) );
  AO21X1 U124 ( .A0(n900), .A1(cnt_data[2]), .B0(n910), .Y(N21) );
  NAND2X1 U125 ( .A(n910), .B(n940), .Y(n920) );
  OAI21XL U126 ( .A0(n910), .A1(n940), .B0(n920), .Y(N22) );
  OR2X1 U127 ( .A(cnt_data[2]), .B(cnt_data[3]), .Y(n950) );
  CLKINVX6 U128 ( .A(rst), .Y(n1030) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_0 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n2), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n3), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n4), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n8), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  INVX1 U1 ( .A(B[0]), .Y(n16) );
  INVX1 U2 ( .A(B[13]), .Y(n3) );
  INVX1 U3 ( .A(B[12]), .Y(n4) );
  INVX1 U4 ( .A(B[3]), .Y(n13) );
  INVX1 U5 ( .A(B[4]), .Y(n12) );
  INVX1 U6 ( .A(B[5]), .Y(n11) );
  INVX1 U7 ( .A(B[6]), .Y(n10) );
  INVX1 U8 ( .A(B[7]), .Y(n9) );
  INVX1 U9 ( .A(B[8]), .Y(n8) );
  INVX1 U10 ( .A(B[9]), .Y(n7) );
  INVX1 U11 ( .A(B[10]), .Y(n6) );
  INVX1 U12 ( .A(B[11]), .Y(n5) );
  INVX1 U13 ( .A(B[2]), .Y(n14) );
  XNOR3X1 U14 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(DIFF[15]) );
  XNOR2XL U15 ( .A(n16), .B(A[0]), .Y(DIFF[0]) );
  NAND2X1 U16 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U17 ( .A(B[1]), .Y(n15) );
  CLKINVX1 U18 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n2) );
endmodule


module FFT_ultrafast2_shift_DW01_add_0 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2XL U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_1 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U2 ( .A(B[15]), .Y(n2) );
  CLKINVX1 U3 ( .A(B[1]), .Y(n16) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U7 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U8 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U9 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U12 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U13 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U14 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U15 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U17 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[14]), .Y(n3) );
  XNOR2X1 U19 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_1 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_2 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n2), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n3), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n4), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n8), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(DIFF[15]) );
  XNOR2X1 U2 ( .A(n16), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n16) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n15) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n14) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n13) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n10) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n9) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n8) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n7) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n5) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n3) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n2) );
endmodule


module FFT_ultrafast2_shift_DW01_add_2 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_3 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n17) );
  NAND2X1 U2 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U3 ( .A(B[1]), .Y(n16) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U5 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U6 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U7 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U8 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U9 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U10 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U11 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U12 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U13 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U14 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U15 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U16 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U17 ( .A(B[14]), .Y(n3) );
  CLKINVX1 U18 ( .A(B[15]), .Y(n2) );
  XNOR2X1 U19 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_3 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_4 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:1] carry;

  ADDFXL U2_13 ( .A(A[13]), .B(n6), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n4), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n16), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n15), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n14), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n13), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n11), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_14 ( .A(A[14]), .B(n7), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n9), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR3X1 U1 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(DIFF[15]) );
  INVX1 U2 ( .A(A[0]), .Y(n1) );
  XNOR2X1 U3 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U4 ( .A(B[0]), .Y(n2) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n8) );
  NAND2X1 U6 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n9) );
  CLKINVX1 U8 ( .A(B[14]), .Y(n7) );
  CLKINVX1 U9 ( .A(B[3]), .Y(n10) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n13) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n14) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n15) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n16) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n3) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n6) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_5 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  XOR3X1 U2_15 ( .A(A[15]), .B(n8), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n7), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n6), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n4), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n17), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n16), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n15), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n14), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n11), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n10), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR2X1 U1 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  NAND2BX1 U2 ( .AN(n2), .B(n1), .Y(carry[1]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n2) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n9) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n10) );
  CLKINVX1 U7 ( .A(B[3]), .Y(n11) );
  CLKINVX1 U8 ( .A(B[14]), .Y(n7) );
  CLKINVX1 U9 ( .A(B[15]), .Y(n8) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n13) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n14) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n15) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n16) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n17) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n3) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n6) );
endmodule


module FFT_ultrafast2_shift_DW01_add_4 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_5 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_6 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  XOR3X1 U2_15 ( .A(A[15]), .B(n8), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n7), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n6), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n4), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n17), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n16), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n15), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n14), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n11), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n10), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND2BX1 U1 ( .AN(n2), .B(n1), .Y(carry[1]) );
  XNOR2X1 U2 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n2) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n9) );
  CLKINVX1 U5 ( .A(B[2]), .Y(n10) );
  CLKINVX1 U6 ( .A(B[3]), .Y(n11) );
  CLKINVX1 U7 ( .A(B[14]), .Y(n7) );
  CLKINVX1 U8 ( .A(B[15]), .Y(n8) );
  CLKINVX1 U9 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n13) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n14) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n15) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n16) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n17) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n3) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n6) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_7 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_13 ( .A(A[13]), .B(n6), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n4), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n17), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n16), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n15), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n14), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n8), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n7), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n10), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n11), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  NAND2BX1 U1 ( .AN(n2), .B(n1), .Y(carry[1]) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  XNOR2X1 U3 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n9) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n10) );
  CLKINVX1 U7 ( .A(B[14]), .Y(n7) );
  CLKINVX1 U8 ( .A(B[15]), .Y(n8) );
  CLKINVX1 U9 ( .A(B[3]), .Y(n11) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n13) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n14) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n15) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n16) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n17) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n3) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n6) );
endmodule


module FFT_ultrafast2_shift_DW01_add_6 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_7 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_12 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n2), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n3), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n4), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n8), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(DIFF[15]) );
  XNOR2X1 U2 ( .A(n16), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n16) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n15) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  INVXL U7 ( .A(B[2]), .Y(n14) );
  INVXL U8 ( .A(B[3]), .Y(n13) );
  INVXL U9 ( .A(B[4]), .Y(n12) );
  INVXL U10 ( .A(B[5]), .Y(n11) );
  INVXL U11 ( .A(B[6]), .Y(n10) );
  INVXL U12 ( .A(B[7]), .Y(n9) );
  INVXL U13 ( .A(B[8]), .Y(n8) );
  INVXL U14 ( .A(B[9]), .Y(n7) );
  INVXL U15 ( .A(B[10]), .Y(n6) );
  INVXL U16 ( .A(B[11]), .Y(n5) );
  INVXL U17 ( .A(B[12]), .Y(n4) );
  INVXL U18 ( .A(B[13]), .Y(n3) );
  INVXL U19 ( .A(B[14]), .Y(n2) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_13 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n2), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n3), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n4), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n8), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(DIFF[15]) );
  XNOR2X1 U2 ( .A(n16), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n16) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n15) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n14) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n13) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n10) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n9) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n8) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n7) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n5) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n3) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n2) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_14 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n2), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n3), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n4), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n7), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n8), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n11), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n12), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n13), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n14), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n15), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(DIFF[15]) );
  XNOR2X1 U2 ( .A(n16), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n16) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n15) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n14) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n13) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n10) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n9) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n8) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n7) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n5) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n3) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n2) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_15 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[15]), .Y(n2) );
  XNOR2X1 U2 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n17) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n16) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n3) );
endmodule


module FFT_ultrafast2_shift_DW01_add_8 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_9 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_10 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_11 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_16 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  XOR3XL U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR2X1 U1 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U3 ( .A(B[1]), .Y(n16) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U6 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U7 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U8 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U9 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U10 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U11 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U12 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U13 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U14 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U15 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U16 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U17 ( .A(B[14]), .Y(n3) );
  CLKINVX1 U18 ( .A(B[15]), .Y(n2) );
  CLKINVX1 U19 ( .A(B[0]), .Y(n17) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_17 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  XNOR2X1 U1 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U2 ( .A(B[14]), .Y(n3) );
  CLKINVX1 U3 ( .A(B[15]), .Y(n2) );
  CLKINVX1 U4 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n16) );
  NAND2X1 U6 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U7 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U8 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U9 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n4) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_18 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  XNOR2X1 U1 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U2 ( .A(B[14]), .Y(n3) );
  CLKINVX1 U3 ( .A(B[15]), .Y(n2) );
  CLKINVX1 U4 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n16) );
  NAND2X1 U6 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U7 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U8 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U9 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n4) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_19 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  XNOR2X1 U1 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U2 ( .A(B[14]), .Y(n3) );
  CLKINVX1 U3 ( .A(B[15]), .Y(n2) );
  CLKINVX1 U4 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U5 ( .A(B[1]), .Y(n16) );
  NAND2X1 U6 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U7 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U8 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U9 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U10 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U12 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U13 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U14 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U15 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U16 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U17 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U18 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U19 ( .A(B[13]), .Y(n4) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_20 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[15]), .Y(n2) );
  XNOR2X1 U2 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n16) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n3) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_21 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[15]), .Y(n2) );
  XNOR2X1 U2 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n16) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n3) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_22 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[15]), .Y(n2) );
  XNOR2X1 U2 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U3 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n16) );
  NAND2X1 U5 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U6 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U7 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U8 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U9 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U10 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U11 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U12 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U13 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U14 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U15 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U16 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U17 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U18 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U19 ( .A(B[14]), .Y(n3) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_23 ( A, B, DIFF );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADDFXL U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .A(A[15]), .B(n2), .C(carry[15]), .Y(DIFF[15]) );
  CLKINVX1 U1 ( .A(B[15]), .Y(n2) );
  CLKINVX1 U2 ( .A(B[0]), .Y(n17) );
  CLKINVX1 U3 ( .A(B[1]), .Y(n16) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n15) );
  CLKINVX1 U7 ( .A(B[3]), .Y(n14) );
  CLKINVX1 U8 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U9 ( .A(B[5]), .Y(n12) );
  CLKINVX1 U10 ( .A(B[6]), .Y(n11) );
  CLKINVX1 U11 ( .A(B[7]), .Y(n10) );
  CLKINVX1 U12 ( .A(B[8]), .Y(n9) );
  CLKINVX1 U13 ( .A(B[9]), .Y(n8) );
  CLKINVX1 U14 ( .A(B[10]), .Y(n7) );
  CLKINVX1 U15 ( .A(B[11]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[12]), .Y(n5) );
  CLKINVX1 U17 ( .A(B[13]), .Y(n4) );
  CLKINVX1 U18 ( .A(B[14]), .Y(n3) );
  XNOR2X1 U19 ( .A(n17), .B(A[0]), .Y(DIFF[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_12 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3XL U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_13 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_14 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_15 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_16 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_17 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_18 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW01_add_19 ( A, B, SUM );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  wire   n1;
  wire   [15:2] carry;

  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module FFT_ultrafast2_shift_DW_mult_uns_8 ( a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        b_31_, b_30_, b_29_, b_28_, b_27_, b_26_, b_25_, b_16_, b_15_, b_14_, 
        b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, 
        b_2_, b_1_, b_0_, product_31_, product_30_, product_29_, product_28_, 
        product_27_, product_26_, product_25_, product_24_, product_23_, 
        product_22_, product_21_, product_20_, product_19_, product_18_, 
        product_17_, product_16_, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_, product_2_, 
        product_1_, product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_, b_31_, b_30_, b_29_, b_28_, b_27_,
         b_26_, b_25_, b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_,
         b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n4, n5, n10, n12, n13, n15, n16, n17, n18, n19, n21, n22, n24,
         n25, n28, n30, n31, n34, n36, n37, n40, n41, n43, n46, n49, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n83, n84, n85, n86, n87, n89, n91, n92, n93, n94, n95, n97, n99,
         n100, n101, n102, n103, n105, n107, n108, n109, n110, n111, n113,
         n115, n116, n117, n118, n119, n121, n123, n124, n125, n126, n127,
         n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n183, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201,
         n203, n204, n205, n206, n207, n209, n211, n212, n213, n214, n216,
         n218, n220, n222, n224, n226, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n239, n240, n241, n243, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n717, n718, n719, n720, n721, n723, n724, n726,
         n727, n728, n729, n730, n731, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n764, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n849, n850, n851, n852, n853;

  XNOR2X1 U694 ( .A(n724), .B(n13), .Y(n670) );
  XNOR2X4 U695 ( .A(n718), .B(n25), .Y(n628) );
  NOR2X2 U696 ( .A(n190), .B(n193), .Y(n188) );
  OAI21X2 U697 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NAND2X1 U698 ( .A(n571), .B(n435), .Y(n214) );
  OAI22X1 U699 ( .A0(n714), .A1(n5), .B0(n713), .B1(n4), .Y(n571) );
  OAI22XL U700 ( .A0(n696), .A1(n12), .B0(n695), .B1(n10), .Y(n553) );
  AOI21X1 U701 ( .A0(n838), .A1(n212), .B0(n209), .Y(n207) );
  OAI22XL U702 ( .A0(n694), .A1(n12), .B0(n693), .B1(n10), .Y(n551) );
  OAI22X1 U703 ( .A0(n658), .A1(n24), .B0(n657), .B1(n21), .Y(n515) );
  CLKBUFX3 U704 ( .A(a_5_), .Y(n13) );
  NOR2X1 U705 ( .A(n388), .B(n395), .Y(n168) );
  ADDFXL U706 ( .A(n377), .B(n559), .CI(n482), .CO(n374), .S(n375) );
  CMPR42X1 U707 ( .A(n497), .B(n381), .C(n382), .D(n373), .ICI(n378), .S(n370), 
        .ICO(n368), .CO(n369) );
  CLKBUFX3 U708 ( .A(n755), .Y(n10) );
  XNOR2X1 U709 ( .A(a_5_), .B(a_6_), .Y(n753) );
  CLKBUFX3 U710 ( .A(a_15_), .Y(n43) );
  AO21X1 U711 ( .A0(n186), .A1(n834), .B0(n183), .Y(n852) );
  OAI22X1 U712 ( .A0(n741), .A1(n573), .B0(n46), .B1(n572), .Y(n246) );
  CLKINVX1 U713 ( .A(n144), .Y(n143) );
  NOR2X1 U714 ( .A(n282), .B(n289), .Y(n117) );
  CLKINVX1 U715 ( .A(n133), .Y(n228) );
  NOR2BXL U716 ( .AN(n49), .B(n750), .Y(n467) );
  XOR2X1 U717 ( .A(a_5_), .B(a_4_), .Y(n738) );
  OR2X1 U718 ( .A(n425), .B(n426), .Y(n833) );
  OR2X1 U719 ( .A(n409), .B(n413), .Y(n834) );
  OR2X1 U720 ( .A(n308), .B(n316), .Y(n835) );
  OR2X1 U721 ( .A(n290), .B(n297), .Y(n836) );
  OR2X1 U722 ( .A(n276), .B(n281), .Y(n837) );
  OR2XL U723 ( .A(n570), .B(n554), .Y(n838) );
  OR2X1 U724 ( .A(n268), .B(n264), .Y(n839) );
  OR2X1 U725 ( .A(n256), .B(n258), .Y(n840) );
  OR2X1 U726 ( .A(n250), .B(n249), .Y(n841) );
  BUFX4 U727 ( .A(n745), .Y(n24) );
  CLKBUFX3 U728 ( .A(n748), .Y(n5) );
  NAND2X2 U729 ( .A(n734), .B(n750), .Y(n742) );
  INVX4 U730 ( .A(n849), .Y(n850) );
  INVX3 U731 ( .A(a_3_), .Y(n849) );
  BUFX4 U732 ( .A(n747), .Y(n12) );
  CLKBUFX3 U733 ( .A(n743), .Y(n36) );
  CLKBUFX3 U734 ( .A(n744), .Y(n30) );
  CMPR42X2 U735 ( .A(n431), .B(n406), .C(n410), .D(n404), .ICI(n407), .S(n402), 
        .ICO(n400), .CO(n401) );
  OAI22X1 U736 ( .A0(n643), .A1(n28), .B0(n30), .B1(n760), .Y(n431) );
  OAI22X1 U737 ( .A0(n697), .A1(n10), .B0(n12), .B1(n849), .Y(n434) );
  OAI22X1 U738 ( .A0(n692), .A1(n10), .B0(n747), .B1(n693), .Y(n550) );
  OAI21X2 U739 ( .A0(n145), .A1(n165), .B0(n146), .Y(n144) );
  XNOR2X2 U740 ( .A(a_3_), .B(a_4_), .Y(n754) );
  XOR2X1 U741 ( .A(n135), .B(n64), .Y(product_18_) );
  CLKINVX1 U742 ( .A(n131), .Y(n129) );
  XNOR2XL U743 ( .A(n37), .B(n731), .Y(n605) );
  XNOR2XL U744 ( .A(n31), .B(n729), .Y(n621) );
  AOI21X2 U745 ( .A0(n132), .A1(n835), .B0(n129), .Y(n127) );
  XNOR2XL U746 ( .A(n727), .B(n13), .Y(n673) );
  XOR2X1 U747 ( .A(n154), .B(n68), .Y(product_14_) );
  CMPR32X2 U748 ( .A(n502), .B(n564), .C(n532), .CO(n410), .S(n411) );
  CLKINVX3 U749 ( .A(n185), .Y(n183) );
  OAI22X1 U750 ( .A0(n690), .A1(n12), .B0(n689), .B1(n755), .Y(n547) );
  XNOR2XL U751 ( .A(n19), .B(n729), .Y(n657) );
  OAI21XL U752 ( .A0(n173), .A1(n171), .B0(n172), .Y(n170) );
  NOR2BX1 U753 ( .AN(n49), .B(n10), .Y(n554) );
  CLKBUFX4 U754 ( .A(a_7_), .Y(n19) );
  OAI21X1 U755 ( .A0(n138), .A1(n142), .B0(n139), .Y(n137) );
  OAI21X2 U756 ( .A0(n127), .A1(n125), .B0(n126), .Y(n124) );
  NAND2XL U757 ( .A(n232), .B(n153), .Y(n68) );
  CLKBUFX2 U758 ( .A(b_4_), .Y(n728) );
  OAI21X2 U759 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  XNOR2XL U760 ( .A(n204), .B(n78), .Y(product_4_) );
  NOR2BXL U761 ( .AN(n49), .B(n28), .Y(n502) );
  NAND2X1 U762 ( .A(n425), .B(n426), .Y(n203) );
  NAND2BXL U763 ( .AN(n49), .B(n1), .Y(n715) );
  INVXL U764 ( .A(n1), .Y(n764) );
  XNOR2XL U765 ( .A(n727), .B(n1), .Y(n709) );
  XNOR2XL U766 ( .A(n728), .B(n1), .Y(n710) );
  XNOR2XL U767 ( .A(n1), .B(n729), .Y(n711) );
  INVX1 U768 ( .A(a_0_), .Y(n756) );
  INVX1 U769 ( .A(n138), .Y(n229) );
  AOI21X1 U770 ( .A0(n164), .A1(n155), .B0(n156), .Y(n154) );
  OAI21XL U771 ( .A0(n154), .A1(n152), .B0(n153), .Y(n151) );
  INVXL U772 ( .A(n149), .Y(n231) );
  NAND2X1 U773 ( .A(n834), .B(n185), .Y(n74) );
  OAI21XL U774 ( .A0(n149), .A1(n153), .B0(n150), .Y(n148) );
  XOR2X1 U775 ( .A(n173), .B(n72), .Y(product_10_) );
  NAND2X1 U776 ( .A(n240), .B(n194), .Y(n76) );
  INVX1 U777 ( .A(n193), .Y(n240) );
  OAI21X1 U778 ( .A0(n207), .A1(n205), .B0(n206), .Y(n204) );
  OAI21XL U779 ( .A0(n87), .A1(n85), .B0(n86), .Y(n84) );
  XOR2XL U780 ( .A(n79), .B(n207), .Y(product_3_) );
  INVXL U781 ( .A(n205), .Y(n243) );
  ADDFX1 U782 ( .A(n547), .B(n531), .CI(n501), .CO(n403), .S(n404) );
  OAI22X1 U783 ( .A0(n642), .A1(n744), .B0(n641), .B1(n28), .Y(n501) );
  OAI22XL U784 ( .A0(n692), .A1(n747), .B0(n691), .B1(n10), .Y(n549) );
  OAI22XL U785 ( .A0(n676), .A1(n17), .B0(n675), .B1(n15), .Y(n533) );
  OAI22XL U786 ( .A0(n622), .A1(n743), .B0(n621), .B1(n34), .Y(n482) );
  OAI22XL U787 ( .A0(n24), .A1(n650), .B0(n649), .B1(n22), .Y(n507) );
  XNOR2X1 U788 ( .A(n730), .B(n1), .Y(n712) );
  XNOR2X1 U789 ( .A(n19), .B(n723), .Y(n651) );
  XNOR2X1 U790 ( .A(n37), .B(n729), .Y(n603) );
  XNOR2X1 U791 ( .A(n724), .B(n850), .Y(n688) );
  XNOR2X1 U792 ( .A(n724), .B(n19), .Y(n652) );
  XNOR2X1 U793 ( .A(n718), .B(n19), .Y(n653) );
  XNOR2X1 U794 ( .A(n726), .B(n19), .Y(n654) );
  XNOR2X1 U795 ( .A(n13), .B(n721), .Y(n667) );
  XNOR2X1 U796 ( .A(n13), .B(b_15_), .Y(n668) );
  OAI22XL U797 ( .A0(n712), .A1(n5), .B0(n711), .B1(n4), .Y(n569) );
  CLKBUFX4 U798 ( .A(a_1_), .Y(n1) );
  OAI21X1 U799 ( .A0(n143), .A1(n141), .B0(n142), .Y(n140) );
  CLKBUFX2 U800 ( .A(b_14_), .Y(n718) );
  INVX3 U801 ( .A(n165), .Y(n164) );
  INVXL U802 ( .A(n174), .Y(n173) );
  CLKBUFX4 U803 ( .A(b_0_), .Y(n49) );
  OAI21X2 U804 ( .A0(n119), .A1(n117), .B0(n118), .Y(n116) );
  OAI21X2 U805 ( .A0(n111), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X2 U806 ( .A0(n103), .A1(n101), .B0(n102), .Y(n100) );
  OAI21X2 U807 ( .A0(n95), .A1(n93), .B0(n94), .Y(n92) );
  INVXL U808 ( .A(n211), .Y(n209) );
  XNOR2X1 U809 ( .A(n851), .B(n69), .Y(product_13_) );
  AO21XL U810 ( .A0(n164), .A1(n234), .B0(n161), .Y(n851) );
  AOI21XL U811 ( .A0(n92), .A1(n841), .B0(n89), .Y(n87) );
  CLKBUFX2 U812 ( .A(b_6_), .Y(n726) );
  CLKBUFX2 U813 ( .A(b_1_), .Y(n731) );
  NOR2X1 U814 ( .A(n350), .B(n360), .Y(n149) );
  INVXL U815 ( .A(n187), .Y(n186) );
  NOR2X1 U816 ( .A(n339), .B(n349), .Y(n141) );
  NOR2X1 U817 ( .A(n328), .B(n338), .Y(n138) );
  NOR2X1 U818 ( .A(n317), .B(n327), .Y(n133) );
  NOR2X1 U819 ( .A(n298), .B(n307), .Y(n125) );
  NAND2XL U820 ( .A(n235), .B(n169), .Y(n71) );
  INVXL U821 ( .A(n168), .Y(n235) );
  NAND2XL U822 ( .A(n236), .B(n172), .Y(n72) );
  XNOR2XL U823 ( .A(n164), .B(n70), .Y(product_12_) );
  NAND2XL U824 ( .A(n234), .B(n163), .Y(n70) );
  INVXL U825 ( .A(n190), .Y(n239) );
  XNOR2X1 U826 ( .A(n852), .B(n73), .Y(product_9_) );
  NOR2X1 U827 ( .A(n370), .B(n379), .Y(n157) );
  NOR2X1 U828 ( .A(n361), .B(n369), .Y(n152) );
  NAND2XL U829 ( .A(n414), .B(n418), .Y(n191) );
  INVXL U830 ( .A(n163), .Y(n161) );
  NOR2X1 U831 ( .A(n275), .B(n269), .Y(n109) );
  NOR2X1 U832 ( .A(n263), .B(n259), .Y(n101) );
  NOR2X1 U833 ( .A(n255), .B(n251), .Y(n93) );
  NOR2X1 U834 ( .A(n248), .B(n247), .Y(n85) );
  ADDHX1 U835 ( .A(n533), .B(n549), .CO(n415), .S(n416) );
  NOR2X1 U836 ( .A(n402), .B(n408), .Y(n179) );
  NOR2BXL U837 ( .AN(n49), .B(n15), .Y(n536) );
  NOR2X1 U838 ( .A(n380), .B(n387), .Y(n162) );
  NOR2BXL U839 ( .AN(n49), .B(n34), .Y(n485) );
  XNOR2XL U840 ( .A(n49), .B(n43), .Y(n588) );
  NOR2X1 U841 ( .A(n396), .B(n401), .Y(n171) );
  NOR2X1 U842 ( .A(n419), .B(n420), .Y(n193) );
  NOR2BXL U843 ( .AN(n49), .B(n46), .Y(n450) );
  NOR2X1 U844 ( .A(n427), .B(n553), .Y(n205) );
  NOR2X1 U845 ( .A(n421), .B(n424), .Y(n197) );
  NAND2BXL U846 ( .AN(n213), .B(n214), .Y(n81) );
  NOR2XL U847 ( .A(n571), .B(n435), .Y(n213) );
  XNOR2XL U848 ( .A(n730), .B(n43), .Y(n586) );
  XNOR2XL U849 ( .A(n731), .B(n43), .Y(n587) );
  NAND2BXL U850 ( .AN(n49), .B(n43), .Y(n589) );
  XNOR2XL U851 ( .A(n727), .B(n43), .Y(n583) );
  XNOR2XL U852 ( .A(n726), .B(n43), .Y(n582) );
  XNOR2XL U853 ( .A(n718), .B(n43), .Y(n581) );
  XNOR2XL U854 ( .A(n724), .B(n43), .Y(n580) );
  XNOR2XL U855 ( .A(n728), .B(n43), .Y(n584) );
  XNOR2XL U856 ( .A(n729), .B(n43), .Y(n585) );
  OAI22XL U857 ( .A0(n24), .A1(n649), .B0(n648), .B1(n22), .Y(n324) );
  OAI22XL U858 ( .A0(n24), .A1(n645), .B0(n644), .B1(n22), .Y(n286) );
  AO21XL U859 ( .A0(n18), .A1(n16), .B0(n662), .Y(n519) );
  AO21XL U860 ( .A0(n5), .A1(n4), .B0(n698), .Y(n555) );
  AO21XL U861 ( .A0(n12), .A1(n10), .B0(n680), .Y(n537) );
  XNOR2XL U862 ( .A(n719), .B(n43), .Y(n575) );
  XNOR2XL U863 ( .A(n718), .B(n43), .Y(n574) );
  XNOR2XL U864 ( .A(n723), .B(n43), .Y(n579) );
  XNOR2XL U865 ( .A(b_15_), .B(n43), .Y(n578) );
  XNOR2XL U866 ( .A(n721), .B(n43), .Y(n577) );
  XNOR2XL U867 ( .A(n43), .B(n720), .Y(n576) );
  AO21XL U868 ( .A0(n30), .A1(n28), .B0(n626), .Y(n486) );
  AO21XL U869 ( .A0(n36), .A1(n34), .B0(n608), .Y(n468) );
  ADDFXL U870 ( .A(n253), .B(n438), .CI(n254), .CO(n250), .S(n251) );
  ADDFXL U871 ( .A(n252), .B(n451), .CI(n437), .CO(n248), .S(n249) );
  AO21XL U872 ( .A0(n742), .A1(n40), .B0(n590), .Y(n451) );
  AO21XL U873 ( .A0(n741), .A1(n46), .B0(n572), .Y(n436) );
  XNOR2XL U874 ( .A(n49), .B(n850), .Y(n696) );
  XNOR2XL U875 ( .A(n850), .B(n731), .Y(n695) );
  XNOR2XL U876 ( .A(b_14_), .B(n13), .Y(n671) );
  XNOR2XL U877 ( .A(n719), .B(n850), .Y(n683) );
  XNOR2XL U878 ( .A(n726), .B(n13), .Y(n672) );
  XNOR2XL U879 ( .A(n726), .B(n25), .Y(n636) );
  XNOR2XL U880 ( .A(n727), .B(n25), .Y(n637) );
  XNOR2XL U881 ( .A(n727), .B(n31), .Y(n619) );
  XNOR2XL U882 ( .A(n727), .B(n19), .Y(n655) );
  XNOR2XL U883 ( .A(n728), .B(n13), .Y(n674) );
  XNOR2XL U884 ( .A(n728), .B(n25), .Y(n638) );
  XNOR2XL U885 ( .A(n730), .B(n19), .Y(n658) );
  XNOR2XL U886 ( .A(n730), .B(n850), .Y(n694) );
  XNOR2XL U887 ( .A(n728), .B(n19), .Y(n656) );
  XNOR2XL U888 ( .A(n728), .B(n31), .Y(n620) );
  XNOR2XL U889 ( .A(n730), .B(n25), .Y(n640) );
  XNOR2XL U890 ( .A(n730), .B(n31), .Y(n622) );
  XNOR2XL U891 ( .A(n730), .B(n37), .Y(n604) );
  XNOR2XL U892 ( .A(n13), .B(n731), .Y(n677) );
  XNOR2XL U893 ( .A(n19), .B(n731), .Y(n659) );
  XNOR2XL U894 ( .A(n850), .B(n729), .Y(n693) );
  CLKBUFX2 U895 ( .A(n753), .Y(n22) );
  CLKBUFX2 U896 ( .A(n753), .Y(n21) );
  XNOR2XL U897 ( .A(n49), .B(n25), .Y(n642) );
  XNOR2XL U898 ( .A(n49), .B(n19), .Y(n660) );
  XNOR2XL U899 ( .A(n49), .B(n13), .Y(n678) );
  XNOR2XL U900 ( .A(n49), .B(n31), .Y(n624) );
  XNOR2XL U901 ( .A(n49), .B(n37), .Y(n606) );
  NAND2BXL U902 ( .AN(n49), .B(n850), .Y(n697) );
  NAND2BXL U903 ( .AN(n49), .B(n19), .Y(n661) );
  NAND2BXL U904 ( .AN(n49), .B(n13), .Y(n679) );
  NAND2BXL U905 ( .AN(n49), .B(n37), .Y(n607) );
  XNOR2XL U906 ( .A(n718), .B(n31), .Y(n617) );
  XNOR2XL U907 ( .A(n724), .B(n25), .Y(n634) );
  XNOR2XL U908 ( .A(n719), .B(n13), .Y(n665) );
  XNOR2XL U909 ( .A(n726), .B(n31), .Y(n618) );
  XNOR2XL U910 ( .A(n727), .B(n37), .Y(n601) );
  XNOR2XL U911 ( .A(n724), .B(n31), .Y(n616) );
  XNOR2XL U912 ( .A(n726), .B(n37), .Y(n600) );
  XNOR2XL U913 ( .A(n718), .B(n850), .Y(n682) );
  XNOR2XL U914 ( .A(n728), .B(n37), .Y(n602) );
  XNOR2XL U915 ( .A(n718), .B(n13), .Y(n664) );
  XNOR2XL U916 ( .A(n19), .B(b_15_), .Y(n650) );
  XNOR2XL U917 ( .A(n31), .B(n731), .Y(n623) );
  XNOR2XL U918 ( .A(n25), .B(n729), .Y(n639) );
  XNOR2XL U919 ( .A(n850), .B(n720), .Y(n684) );
  XNOR2XL U920 ( .A(n13), .B(n720), .Y(n666) );
  NAND2BXL U921 ( .AN(n49), .B(n31), .Y(n625) );
  XNOR2XL U922 ( .A(n719), .B(n19), .Y(n647) );
  XNOR2XL U923 ( .A(n718), .B(n37), .Y(n599) );
  XNOR2XL U924 ( .A(n724), .B(n37), .Y(n598) );
  XNOR2XL U925 ( .A(n719), .B(n25), .Y(n629) );
  XNOR2XL U926 ( .A(n719), .B(n31), .Y(n611) );
  XNOR2XL U927 ( .A(n718), .B(n19), .Y(n646) );
  XNOR2XL U928 ( .A(n718), .B(n31), .Y(n610) );
  XNOR2XL U929 ( .A(n850), .B(n717), .Y(n681) );
  XNOR2XL U930 ( .A(n25), .B(n717), .Y(n632) );
  XNOR2XL U931 ( .A(n31), .B(n717), .Y(n614) );
  XNOR2XL U932 ( .A(n13), .B(n717), .Y(n663) );
  XNOR2XL U933 ( .A(n37), .B(b_15_), .Y(n596) );
  XNOR2XL U934 ( .A(n25), .B(n723), .Y(n633) );
  XNOR2XL U935 ( .A(n31), .B(n723), .Y(n615) );
  XNOR2XL U936 ( .A(n37), .B(n723), .Y(n597) );
  XNOR2XL U937 ( .A(n25), .B(n721), .Y(n631) );
  XNOR2XL U938 ( .A(n31), .B(n721), .Y(n613) );
  XNOR2XL U939 ( .A(n37), .B(n721), .Y(n595) );
  XNOR2XL U940 ( .A(n25), .B(n720), .Y(n630) );
  XNOR2XL U941 ( .A(n31), .B(n720), .Y(n612) );
  XNOR2XL U942 ( .A(n850), .B(b_31_), .Y(n680) );
  XNOR2XL U943 ( .A(n13), .B(b_30_), .Y(n662) );
  XNOR2XL U944 ( .A(n719), .B(n37), .Y(n593) );
  XNOR2XL U945 ( .A(n718), .B(n37), .Y(n592) );
  XNOR2XL U946 ( .A(n25), .B(n717), .Y(n627) );
  XNOR2XL U947 ( .A(n37), .B(n720), .Y(n594) );
  XNOR2XL U948 ( .A(n25), .B(b_28_), .Y(n626) );
  XNOR2XL U949 ( .A(n31), .B(n717), .Y(n609) );
  XNOR2XL U950 ( .A(n37), .B(n717), .Y(n591) );
  XNOR2XL U951 ( .A(n31), .B(b_27_), .Y(n608) );
  XNOR2XL U952 ( .A(n37), .B(b_26_), .Y(n590) );
  XNOR2X1 U953 ( .A(a_1_), .B(a_2_), .Y(n755) );
  XNOR2X1 U954 ( .A(a_7_), .B(a_8_), .Y(n752) );
  XNOR2X1 U955 ( .A(a_11_), .B(a_12_), .Y(n750) );
  XNOR2X1 U956 ( .A(a_9_), .B(a_10_), .Y(n751) );
  CLKBUFX3 U957 ( .A(a_9_), .Y(n25) );
  NAND2X4 U958 ( .A(n738), .B(n754), .Y(n746) );
  CLKBUFX3 U959 ( .A(a_11_), .Y(n31) );
  CLKBUFX3 U960 ( .A(a_13_), .Y(n37) );
  XNOR2X1 U961 ( .A(a_13_), .B(a_14_), .Y(n749) );
  NAND2X4 U962 ( .A(n749), .B(n733), .Y(n741) );
  XNOR2X1 U963 ( .A(n140), .B(n65), .Y(product_17_) );
  NAND2X1 U964 ( .A(n229), .B(n139), .Y(n65) );
  XNOR2X1 U965 ( .A(n132), .B(n63), .Y(product_19_) );
  NAND2X1 U966 ( .A(n835), .B(n131), .Y(n63) );
  AOI21X1 U967 ( .A0(n144), .A1(n136), .B0(n137), .Y(n135) );
  NOR2X1 U968 ( .A(n141), .B(n138), .Y(n136) );
  OAI21X1 U969 ( .A0(n135), .A1(n133), .B0(n134), .Y(n132) );
  XOR2X1 U970 ( .A(n127), .B(n62), .Y(product_20_) );
  NAND2X1 U971 ( .A(n226), .B(n126), .Y(n62) );
  CLKINVX1 U972 ( .A(n125), .Y(n226) );
  NAND2X1 U973 ( .A(n228), .B(n134), .Y(n64) );
  XOR2X1 U974 ( .A(n143), .B(n66), .Y(product_16_) );
  NAND2X1 U975 ( .A(n230), .B(n142), .Y(n66) );
  CLKINVX1 U976 ( .A(n141), .Y(n230) );
  XNOR2X1 U977 ( .A(n80), .B(n212), .Y(product_2_) );
  NAND2X1 U978 ( .A(n838), .B(n211), .Y(n80) );
  XNOR2X1 U979 ( .A(n186), .B(n74), .Y(product_8_) );
  XNOR2X1 U980 ( .A(n151), .B(n67), .Y(product_15_) );
  NAND2X1 U981 ( .A(n231), .B(n150), .Y(n67) );
  XNOR2X1 U982 ( .A(n92), .B(n53), .Y(product_29_) );
  NAND2X1 U983 ( .A(n841), .B(n91), .Y(n53) );
  XNOR2X1 U984 ( .A(n100), .B(n55), .Y(product_27_) );
  NAND2X1 U985 ( .A(n840), .B(n99), .Y(n55) );
  XNOR2X1 U986 ( .A(n108), .B(n57), .Y(product_25_) );
  NAND2X1 U987 ( .A(n839), .B(n107), .Y(n57) );
  XNOR2X1 U988 ( .A(n116), .B(n59), .Y(product_23_) );
  NAND2X1 U989 ( .A(n837), .B(n115), .Y(n59) );
  XNOR2X1 U990 ( .A(n124), .B(n61), .Y(product_21_) );
  NAND2X1 U991 ( .A(n836), .B(n123), .Y(n61) );
  NAND2X1 U992 ( .A(n147), .B(n155), .Y(n145) );
  AOI21X1 U993 ( .A0(n156), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U994 ( .A(n152), .B(n149), .Y(n147) );
  AOI21X1 U995 ( .A0(n124), .A1(n836), .B0(n121), .Y(n119) );
  CLKINVX1 U996 ( .A(n123), .Y(n121) );
  AOI21X1 U997 ( .A0(n116), .A1(n837), .B0(n113), .Y(n111) );
  CLKINVX1 U998 ( .A(n115), .Y(n113) );
  AOI21X1 U999 ( .A0(n108), .A1(n839), .B0(n105), .Y(n103) );
  CLKINVX1 U1000 ( .A(n107), .Y(n105) );
  AOI21X1 U1001 ( .A0(n100), .A1(n840), .B0(n97), .Y(n95) );
  CLKINVX1 U1002 ( .A(n99), .Y(n97) );
  CLKINVX1 U1003 ( .A(n91), .Y(n89) );
  CLKBUFX3 U1004 ( .A(b_15_), .Y(n717) );
  CLKBUFX3 U1005 ( .A(b_11_), .Y(n721) );
  CLKBUFX3 U1006 ( .A(b_5_), .Y(n727) );
  CLKBUFX3 U1007 ( .A(b_13_), .Y(n719) );
  CLKBUFX3 U1008 ( .A(b_2_), .Y(n730) );
  CLKBUFX3 U1009 ( .A(b_8_), .Y(n724) );
  NAND2X1 U1010 ( .A(n339), .B(n349), .Y(n142) );
  NAND2X1 U1011 ( .A(n308), .B(n316), .Y(n131) );
  NAND2X1 U1012 ( .A(n350), .B(n360), .Y(n150) );
  NAND2X1 U1013 ( .A(n328), .B(n338), .Y(n139) );
  NAND2X1 U1014 ( .A(n317), .B(n327), .Y(n134) );
  NAND2X1 U1015 ( .A(n233), .B(n158), .Y(n69) );
  CLKINVX1 U1016 ( .A(n157), .Y(n233) );
  XOR2X1 U1017 ( .A(n87), .B(n52), .Y(product_30_) );
  NAND2X1 U1018 ( .A(n216), .B(n86), .Y(n52) );
  CLKINVX1 U1019 ( .A(n85), .Y(n216) );
  XOR2X1 U1020 ( .A(n95), .B(n54), .Y(product_28_) );
  NAND2X1 U1021 ( .A(n218), .B(n94), .Y(n54) );
  CLKINVX1 U1022 ( .A(n93), .Y(n218) );
  XOR2X1 U1023 ( .A(n103), .B(n56), .Y(product_26_) );
  NAND2X1 U1024 ( .A(n220), .B(n102), .Y(n56) );
  CLKINVX1 U1025 ( .A(n101), .Y(n220) );
  XOR2X1 U1026 ( .A(n111), .B(n58), .Y(product_24_) );
  NAND2X1 U1027 ( .A(n222), .B(n110), .Y(n58) );
  CLKINVX1 U1028 ( .A(n109), .Y(n222) );
  XOR2X1 U1029 ( .A(n119), .B(n60), .Y(product_22_) );
  NAND2X1 U1030 ( .A(n224), .B(n118), .Y(n60) );
  CLKINVX1 U1031 ( .A(n117), .Y(n224) );
  CLKINVX1 U1032 ( .A(n152), .Y(n232) );
  CLKINVX1 U1033 ( .A(n196), .Y(n195) );
  NAND2X1 U1034 ( .A(n298), .B(n307), .Y(n126) );
  NAND2X1 U1035 ( .A(n833), .B(n203), .Y(n78) );
  XNOR2X1 U1036 ( .A(n170), .B(n71), .Y(product_11_) );
  XNOR2X1 U1037 ( .A(n84), .B(n51), .Y(product_31_) );
  NAND2X1 U1038 ( .A(n853), .B(n83), .Y(n51) );
  NAND2X1 U1039 ( .A(n436), .B(n246), .Y(n83) );
  CLKINVX1 U1040 ( .A(n162), .Y(n234) );
  CMPR42X1 U1041 ( .A(n344), .B(n334), .C(n341), .D(n331), .ICI(n337), .S(n328), .ICO(n326), .CO(n327) );
  CMPR42X1 U1042 ( .A(n366), .B(n356), .C(n363), .D(n353), .ICI(n359), .S(n350), .ICO(n348), .CO(n349) );
  CMPR42X1 U1043 ( .A(n374), .B(n367), .C(n372), .D(n364), .ICI(n368), .S(n361), .ICO(n359), .CO(n360) );
  CMPR42X1 U1044 ( .A(n345), .B(n355), .C(n352), .D(n342), .ICI(n348), .S(n339), .ICO(n337), .CO(n338) );
  CMPR42X1 U1045 ( .A(n318), .B(n314), .C(n311), .D(n319), .ICI(n315), .S(n308), .ICO(n306), .CO(n307) );
  CMPR42X1 U1046 ( .A(n329), .B(n333), .C(n330), .D(n320), .ICI(n326), .S(n317), .ICO(n315), .CO(n316) );
  CMPR42X1 U1047 ( .A(n303), .B(n309), .C(n310), .D(n301), .ICI(n306), .S(n298), .ICO(n296), .CO(n297) );
  AOI21X1 U1048 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U1049 ( .A0(n187), .A1(n175), .B0(n176), .Y(n174) );
  NAND2X1 U1050 ( .A(n177), .B(n834), .Y(n175) );
  AOI21X1 U1051 ( .A0(n177), .A1(n183), .B0(n178), .Y(n176) );
  CLKINVX1 U1052 ( .A(n179), .Y(n177) );
  AOI21X1 U1053 ( .A0(n174), .A1(n166), .B0(n167), .Y(n165) );
  NOR2X1 U1054 ( .A(n168), .B(n171), .Y(n166) );
  OAI21XL U1055 ( .A0(n168), .A1(n172), .B0(n169), .Y(n167) );
  NOR2X1 U1056 ( .A(n414), .B(n418), .Y(n190) );
  AOI21X1 U1057 ( .A0(n204), .A1(n833), .B0(n201), .Y(n199) );
  CLKINVX1 U1058 ( .A(n203), .Y(n201) );
  OAI21X1 U1059 ( .A0(n157), .A1(n163), .B0(n158), .Y(n156) );
  XNOR2X1 U1060 ( .A(n192), .B(n75), .Y(product_7_) );
  NAND2X1 U1061 ( .A(n239), .B(n191), .Y(n75) );
  OAI21XL U1062 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2X1 U1063 ( .A(n361), .B(n369), .Y(n153) );
  NOR2X1 U1064 ( .A(n157), .B(n162), .Y(n155) );
  NAND2X1 U1065 ( .A(n570), .B(n554), .Y(n211) );
  NAND2X1 U1066 ( .A(n409), .B(n413), .Y(n185) );
  NAND2X1 U1067 ( .A(n370), .B(n379), .Y(n158) );
  NAND2X1 U1068 ( .A(n177), .B(n180), .Y(n73) );
  NAND2X1 U1069 ( .A(n243), .B(n206), .Y(n79) );
  XOR2X1 U1070 ( .A(n195), .B(n76), .Y(product_6_) );
  CLKINVX1 U1071 ( .A(n171), .Y(n236) );
  XOR2X1 U1072 ( .A(n199), .B(n77), .Y(product_5_) );
  NAND2X1 U1073 ( .A(n241), .B(n198), .Y(n77) );
  CLKINVX1 U1074 ( .A(n197), .Y(n241) );
  CLKINVX1 U1075 ( .A(n214), .Y(n212) );
  CLKINVX1 U1076 ( .A(n324), .Y(n325) );
  CLKINVX1 U1077 ( .A(n180), .Y(n178) );
  NAND2X1 U1078 ( .A(n268), .B(n264), .Y(n107) );
  NAND2X1 U1079 ( .A(n290), .B(n297), .Y(n123) );
  NAND2X1 U1080 ( .A(n276), .B(n281), .Y(n115) );
  NAND2X1 U1081 ( .A(n275), .B(n269), .Y(n110) );
  NAND2X1 U1082 ( .A(n282), .B(n289), .Y(n118) );
  CLKINVX1 U1083 ( .A(n286), .Y(n287) );
  NAND2X1 U1084 ( .A(n256), .B(n258), .Y(n99) );
  NAND2X1 U1085 ( .A(n263), .B(n259), .Y(n102) );
  NAND2X1 U1086 ( .A(n250), .B(n249), .Y(n91) );
  NAND2X1 U1087 ( .A(n255), .B(n251), .Y(n94) );
  NAND2X1 U1088 ( .A(n248), .B(n247), .Y(n86) );
  CLKINVX1 U1089 ( .A(n246), .Y(n247) );
  OR2X1 U1090 ( .A(n436), .B(n246), .Y(n853) );
  OAI22X1 U1091 ( .A0(n712), .A1(n4), .B0(n5), .B1(n713), .Y(n570) );
  CMPR42X1 U1092 ( .A(n518), .B(n550), .C(n534), .D(n566), .ICI(n422), .S(n419), .ICO(n417), .CO(n418) );
  OAI22XL U1093 ( .A0(n709), .A1(n5), .B0(n708), .B1(n4), .Y(n566) );
  OAI22XL U1094 ( .A0(n676), .A1(n15), .B0(n17), .B1(n677), .Y(n534) );
  NOR2BX1 U1095 ( .AN(n49), .B(n21), .Y(n518) );
  CMPR42X1 U1096 ( .A(n516), .B(n548), .C(n415), .D(n411), .ICI(n412), .S(n409), .ICO(n407), .CO(n408) );
  OAI22XL U1097 ( .A0(n691), .A1(n747), .B0(n690), .B1(n10), .Y(n548) );
  OAI22XL U1098 ( .A0(n658), .A1(n21), .B0(n24), .B1(n659), .Y(n516) );
  CMPR42X1 U1099 ( .A(n565), .B(n432), .C(n517), .D(n416), .ICI(n417), .S(n414), .ICO(n412), .CO(n413) );
  OAI22XL U1100 ( .A0(n661), .A1(n22), .B0(n24), .B1(n761), .Y(n432) );
  OAI22XL U1101 ( .A0(n660), .A1(n24), .B0(n659), .B1(n21), .Y(n517) );
  OAI22XL U1102 ( .A0(n708), .A1(n5), .B0(n707), .B1(n4), .Y(n565) );
  OAI22XL U1103 ( .A0(n638), .A1(n30), .B0(n637), .B1(n28), .Y(n497) );
  CMPR42X1 U1104 ( .A(n528), .B(n385), .C(n390), .D(n383), .ICI(n386), .S(n380), .ICO(n378), .CO(n379) );
  OAI22XL U1105 ( .A0(n671), .A1(n17), .B0(n670), .B1(n15), .Y(n528) );
  CLKBUFX3 U1106 ( .A(b_12_), .Y(n720) );
  CLKBUFX3 U1107 ( .A(b_3_), .Y(n729) );
  CLKBUFX3 U1108 ( .A(b_9_), .Y(n723) );
  OAI22XL U1109 ( .A0(n638), .A1(n28), .B0(n744), .B1(n639), .Y(n498) );
  OAI22XL U1110 ( .A0(n700), .A1(n5), .B0(n699), .B1(n4), .Y(n557) );
  OAI22XL U1111 ( .A0(n700), .A1(n4), .B0(n701), .B1(n5), .Y(n558) );
  OAI22XL U1112 ( .A0(n682), .A1(n12), .B0(n681), .B1(n10), .Y(n539) );
  OAI22XL U1113 ( .A0(n30), .A1(n633), .B0(n632), .B1(n28), .Y(n492) );
  OAI22XL U1114 ( .A0(n689), .A1(n12), .B0(n688), .B1(n10), .Y(n546) );
  ADDFX2 U1115 ( .A(n536), .B(n568), .CI(n552), .CO(n424), .S(n425) );
  OAI22XL U1116 ( .A0(n694), .A1(n10), .B0(n747), .B1(n695), .Y(n552) );
  OAI22XL U1117 ( .A0(n710), .A1(n4), .B0(n5), .B1(n711), .Y(n568) );
  ADDHXL U1118 ( .A(n563), .B(n515), .CO(n405), .S(n406) );
  OAI22XL U1119 ( .A0(n706), .A1(n5), .B0(n705), .B1(n4), .Y(n563) );
  ADDHXL U1120 ( .A(n524), .B(n556), .CO(n346), .S(n347) );
  OAI22XL U1121 ( .A0(n5), .A1(n699), .B0(n698), .B1(n4), .Y(n556) );
  OAI22XL U1122 ( .A0(n18), .A1(n667), .B0(n666), .B1(n16), .Y(n524) );
  ADDHXL U1123 ( .A(n561), .B(n545), .CO(n392), .S(n393) );
  OAI22XL U1124 ( .A0(n5), .A1(n704), .B0(n703), .B1(n4), .Y(n561) );
  OAI22XL U1125 ( .A0(n688), .A1(n747), .B0(n687), .B1(n10), .Y(n545) );
  ADDHXL U1126 ( .A(n525), .B(n509), .CO(n357), .S(n358) );
  OAI22XL U1127 ( .A0(n18), .A1(n668), .B0(n667), .B1(n16), .Y(n525) );
  OAI22XL U1128 ( .A0(n652), .A1(n24), .B0(n651), .B1(n22), .Y(n509) );
  NAND2X1 U1129 ( .A(n380), .B(n387), .Y(n163) );
  NAND2X1 U1130 ( .A(n396), .B(n401), .Y(n172) );
  CMPR42X1 U1131 ( .A(n358), .B(n541), .C(n464), .D(n449), .ICI(n362), .S(n356), .ICO(n354), .CO(n355) );
  OAI22XL U1132 ( .A0(n683), .A1(n10), .B0(n12), .B1(n684), .Y(n541) );
  OAI22XL U1133 ( .A0(n588), .A1(n741), .B0(n46), .B1(n587), .Y(n449) );
  OAI22XL U1134 ( .A0(n604), .A1(n41), .B0(n603), .B1(n40), .Y(n464) );
  CMPR42X1 U1135 ( .A(n491), .B(n324), .C(n537), .D(n476), .ICI(n445), .S(n314), .ICO(n312), .CO(n313) );
  OAI22XL U1136 ( .A0(n616), .A1(n36), .B0(n615), .B1(n34), .Y(n476) );
  OAI22XL U1137 ( .A0(n584), .A1(n741), .B0(n583), .B1(n46), .Y(n445) );
  CMPR42X1 U1138 ( .A(n493), .B(n346), .C(n523), .D(n336), .ICI(n343), .S(n334), .ICO(n332), .CO(n333) );
  OAI22XL U1139 ( .A0(n634), .A1(n30), .B0(n633), .B1(n28), .Y(n493) );
  OAI22XL U1140 ( .A0(n665), .A1(n16), .B0(n18), .B1(n666), .Y(n523) );
  XNOR2X1 U1141 ( .A(n555), .B(n507), .Y(n336) );
  CMPR42X1 U1142 ( .A(n542), .B(n526), .C(n376), .D(n450), .ICI(n496), .S(n367), .ICO(n365), .CO(n366) );
  OAI22XL U1143 ( .A0(n637), .A1(n30), .B0(n636), .B1(n28), .Y(n496) );
  OAI22XL U1144 ( .A0(n18), .A1(n669), .B0(n668), .B1(n16), .Y(n526) );
  OAI22XL U1145 ( .A0(n12), .A1(n685), .B0(n684), .B1(n10), .Y(n542) );
  NAND2X1 U1146 ( .A(n419), .B(n420), .Y(n194) );
  CMPR42X1 U1147 ( .A(n508), .B(n347), .C(n357), .D(n540), .ICI(n479), .S(n345), .ICO(n343), .CO(n344) );
  OAI22XL U1148 ( .A0(n619), .A1(n743), .B0(n618), .B1(n34), .Y(n479) );
  OAI22XL U1149 ( .A0(n24), .A1(n651), .B0(n650), .B1(n22), .Y(n508) );
  OAI22XL U1150 ( .A0(n682), .A1(n10), .B0(n683), .B1(n12), .Y(n540) );
  NAND2X1 U1151 ( .A(n402), .B(n408), .Y(n180) );
  CMPR42X1 U1152 ( .A(n506), .B(n321), .C(n521), .D(n460), .ICI(n322), .S(n311), .ICO(n309), .CO(n310) );
  OAI22XL U1153 ( .A0(n600), .A1(n41), .B0(n599), .B1(n40), .Y(n460) );
  OAI22XL U1154 ( .A0(n664), .A1(n18), .B0(n663), .B1(n16), .Y(n521) );
  OAI22XL U1155 ( .A0(n647), .A1(n22), .B0(n24), .B1(n648), .Y(n506) );
  CMPR42X1 U1156 ( .A(n500), .B(n405), .C(n403), .D(n400), .ICI(n399), .S(n396), .ICO(n394), .CO(n395) );
  OAI22XL U1157 ( .A0(n640), .A1(n28), .B0(n744), .B1(n641), .Y(n500) );
  CMPR42X1 U1158 ( .A(n393), .B(n499), .C(n529), .D(n484), .ICI(n397), .S(n391), .ICO(n389), .CO(n390) );
  OAI22XL U1159 ( .A0(n624), .A1(n36), .B0(n623), .B1(n34), .Y(n484) );
  OAI22XL U1160 ( .A0(n672), .A1(n17), .B0(n671), .B1(n15), .Y(n529) );
  OAI22XL U1161 ( .A0(n640), .A1(n744), .B0(n639), .B1(n28), .Y(n499) );
  CMPR42X1 U1162 ( .A(n467), .B(n498), .C(n483), .D(n512), .ICI(n389), .S(n383), .ICO(n381), .CO(n382) );
  OAI22XL U1163 ( .A0(n655), .A1(n24), .B0(n654), .B1(n21), .Y(n512) );
  OAI22XL U1164 ( .A0(n622), .A1(n34), .B0(n743), .B1(n623), .Y(n483) );
  CMPR42X1 U1165 ( .A(n494), .B(n463), .C(n448), .D(n354), .ICI(n351), .S(n342), .ICO(n340), .CO(n341) );
  OAI22XL U1166 ( .A0(n586), .A1(n46), .B0(n741), .B1(n587), .Y(n448) );
  OAI22XL U1167 ( .A0(n602), .A1(n40), .B0(n41), .B1(n603), .Y(n463) );
  OAI22XL U1168 ( .A0(n628), .A1(n30), .B0(n634), .B1(n28), .Y(n494) );
  CMPR42X1 U1169 ( .A(n558), .B(n510), .C(n481), .D(n465), .ICI(n371), .S(n364), .ICO(n362), .CO(n363) );
  OAI22XL U1170 ( .A0(n604), .A1(n750), .B0(n41), .B1(n605), .Y(n465) );
  OAI22XL U1171 ( .A0(n620), .A1(n34), .B0(n36), .B1(n621), .Y(n481) );
  OAI22XL U1172 ( .A0(n653), .A1(n24), .B0(n652), .B1(n21), .Y(n510) );
  NAND2X1 U1173 ( .A(n388), .B(n395), .Y(n169) );
  CMPR42X1 U1174 ( .A(n511), .B(n429), .C(n466), .D(n384), .ICI(n375), .S(n373), .ICO(n371), .CO(n372) );
  OAI22XL U1175 ( .A0(n607), .A1(n40), .B0(n742), .B1(n758), .Y(n429) );
  OAI22XL U1176 ( .A0(n606), .A1(n41), .B0(n605), .B1(n750), .Y(n466) );
  OAI22XL U1177 ( .A0(n654), .A1(n24), .B0(n653), .B1(n21), .Y(n511) );
  CMPR42X1 U1178 ( .A(n557), .B(n495), .C(n480), .D(n428), .ICI(n365), .S(n353), .ICO(n351), .CO(n352) );
  OAI22XL U1179 ( .A0(n589), .A1(n46), .B0(n741), .B1(n757), .Y(n428) );
  OAI22XL U1180 ( .A0(n620), .A1(n743), .B0(n619), .B1(n34), .Y(n480) );
  OAI22XL U1181 ( .A0(n636), .A1(n744), .B0(n628), .B1(n28), .Y(n495) );
  CMPR42X1 U1182 ( .A(n539), .B(n447), .C(n478), .D(n462), .ICI(n340), .S(n331), .ICO(n329), .CO(n330) );
  OAI22XL U1183 ( .A0(n602), .A1(n41), .B0(n601), .B1(n40), .Y(n462) );
  OAI22XL U1184 ( .A0(n618), .A1(n743), .B0(n617), .B1(n34), .Y(n478) );
  OAI22XL U1185 ( .A0(n586), .A1(n741), .B0(n46), .B1(n585), .Y(n447) );
  CMPR42X1 U1186 ( .A(n522), .B(n477), .C(n446), .D(n332), .ICI(n323), .S(n320), .ICO(n318), .CO(n319) );
  OAI22XL U1187 ( .A0(n584), .A1(n749), .B0(n741), .B1(n585), .Y(n446) );
  OAI22XL U1188 ( .A0(n617), .A1(n743), .B0(n616), .B1(n34), .Y(n477) );
  OAI22XL U1189 ( .A0(n664), .A1(n16), .B0(n665), .B1(n18), .Y(n522) );
  CMPR42X1 U1190 ( .A(n312), .B(n505), .C(n459), .D(n444), .ICI(n313), .S(n301), .ICO(n299), .CO(n300) );
  OAI22XL U1191 ( .A0(n583), .A1(n741), .B0(n582), .B1(n749), .Y(n444) );
  OAI22XL U1192 ( .A0(n599), .A1(n41), .B0(n598), .B1(n40), .Y(n459) );
  OAI22XL U1193 ( .A0(n646), .A1(n22), .B0(n647), .B1(n24), .Y(n505) );
  CLKINVX1 U1194 ( .A(n81), .Y(product_1_) );
  NAND2X1 U1195 ( .A(n427), .B(n553), .Y(n206) );
  CMPR42X1 U1196 ( .A(n562), .B(n485), .C(n546), .D(n514), .ICI(n530), .S(n399), .ICO(n397), .CO(n398) );
  OAI22XL U1197 ( .A0(n673), .A1(n17), .B0(n672), .B1(n15), .Y(n530) );
  OAI22XL U1198 ( .A0(n5), .A1(n705), .B0(n704), .B1(n4), .Y(n562) );
  OAI22XL U1199 ( .A0(n656), .A1(n21), .B0(n24), .B1(n657), .Y(n514) );
  NAND2X1 U1200 ( .A(n421), .B(n424), .Y(n198) );
  CMPR42X1 U1201 ( .A(n492), .B(n538), .C(n325), .D(n335), .ICI(n461), .S(n323), .ICO(n321), .CO(n322) );
  OAI22XL U1202 ( .A0(n601), .A1(n41), .B0(n600), .B1(n40), .Y(n461) );
  OAI22XL U1203 ( .A0(n12), .A1(n681), .B0(n680), .B1(n10), .Y(n538) );
  OR2X1 U1204 ( .A(n555), .B(n507), .Y(n335) );
  ADDHXL U1205 ( .A(n543), .B(n527), .CO(n376), .S(n377) );
  OAI22XL U1206 ( .A0(n12), .A1(n686), .B0(n685), .B1(n10), .Y(n543) );
  OAI22XL U1207 ( .A0(n670), .A1(n17), .B0(n669), .B1(n16), .Y(n527) );
  OAI22XL U1208 ( .A0(n674), .A1(n15), .B0(n17), .B1(n675), .Y(n532) );
  OAI22XL U1209 ( .A0(n707), .A1(n5), .B0(n706), .B1(n4), .Y(n564) );
  OAI22XL U1210 ( .A0(n674), .A1(n17), .B0(n673), .B1(n15), .Y(n531) );
  ADDFXL U1211 ( .A(n544), .B(n560), .CI(n392), .CO(n384), .S(n385) );
  OAI22XL U1212 ( .A0(n5), .A1(n703), .B0(n702), .B1(n4), .Y(n560) );
  OAI22XL U1213 ( .A0(n12), .A1(n687), .B0(n686), .B1(n10), .Y(n544) );
  ADDHXL U1214 ( .A(n551), .B(n567), .CO(n422), .S(n423) );
  OAI22XL U1215 ( .A0(n710), .A1(n5), .B0(n709), .B1(n4), .Y(n567) );
  OAI22XL U1216 ( .A0(n701), .A1(n4), .B0(n5), .B1(n702), .Y(n559) );
  OAI22XL U1217 ( .A0(n30), .A1(n631), .B0(n630), .B1(n28), .Y(n304) );
  OAI22XL U1218 ( .A0(n741), .A1(n579), .B0(n46), .B1(n578), .Y(n272) );
  CMPR42X1 U1219 ( .A(n504), .B(n299), .C(n293), .D(n300), .ICI(n296), .S(n290), .ICO(n288), .CO(n289) );
  OAI22XL U1220 ( .A0(n646), .A1(n24), .B0(n645), .B1(n22), .Y(n504) );
  CMPR42X1 U1221 ( .A(n472), .B(n283), .C(n279), .D(n284), .ICI(n280), .S(n276), .ICO(n274), .CO(n275) );
  OAI22XL U1222 ( .A0(n611), .A1(n34), .B0(n36), .B1(n612), .Y(n472) );
  CMPR42X1 U1223 ( .A(n489), .B(n291), .C(n285), .D(n292), .ICI(n288), .S(n282), .ICO(n280), .CO(n281) );
  OAI22XL U1224 ( .A0(n628), .A1(n28), .B0(n629), .B1(n30), .Y(n489) );
  CMPR42X1 U1225 ( .A(n454), .B(n270), .C(n266), .D(n470), .ICI(n267), .S(n264), .ICO(n262), .CO(n263) );
  OAI22XL U1226 ( .A0(n610), .A1(n36), .B0(n609), .B1(n34), .Y(n470) );
  OAI22XL U1227 ( .A0(n593), .A1(n40), .B0(n742), .B1(n594), .Y(n454) );
  CMPR42X1 U1228 ( .A(n277), .B(n271), .C(n471), .D(n278), .ICI(n274), .S(n269), .ICO(n267), .CO(n268) );
  OAI22XL U1229 ( .A0(n610), .A1(n34), .B0(n611), .B1(n36), .Y(n471) );
  OAI22XL U1230 ( .A0(n742), .A1(n596), .B0(n595), .B1(n40), .Y(n456) );
  OAI22XL U1231 ( .A0(n30), .A1(n632), .B0(n631), .B1(n28), .Y(n491) );
  CMPR42X1 U1232 ( .A(n458), .B(n490), .C(n302), .D(n295), .ICI(n443), .S(n293), .ICO(n291), .CO(n292) );
  OAI22XL U1233 ( .A0(n582), .A1(n741), .B0(n581), .B1(n749), .Y(n443) );
  OAI22XL U1234 ( .A0(n598), .A1(n41), .B0(n597), .B1(n40), .Y(n458) );
  OAI22XL U1235 ( .A0(n629), .A1(n28), .B0(n30), .B1(n630), .Y(n490) );
  CMPR42X1 U1236 ( .A(n286), .B(n456), .C(n503), .D(n441), .ICI(n488), .S(n279), .ICO(n277), .CO(n278) );
  OAI22XL U1237 ( .A0(n628), .A1(n30), .B0(n627), .B1(n28), .Y(n488) );
  OAI22XL U1238 ( .A0(n580), .A1(n741), .B0(n46), .B1(n579), .Y(n441) );
  AO21X1 U1239 ( .A0(n24), .A1(n22), .B0(n644), .Y(n503) );
  CMPR42X1 U1240 ( .A(n457), .B(n473), .C(n287), .D(n294), .ICI(n442), .S(n285), .ICO(n283), .CO(n284) );
  OAI22XL U1241 ( .A0(n581), .A1(n741), .B0(n580), .B1(n46), .Y(n442) );
  OAI22XL U1242 ( .A0(n36), .A1(n613), .B0(n612), .B1(n34), .Y(n473) );
  OAI22XL U1243 ( .A0(n742), .A1(n597), .B0(n596), .B1(n40), .Y(n457) );
  NOR2BX1 U1244 ( .AN(n49), .B(n4), .Y(product_0_) );
  ADDFXL U1245 ( .A(n455), .B(n487), .CI(n273), .CO(n270), .S(n271) );
  OAI22XL U1246 ( .A0(n742), .A1(n595), .B0(n594), .B1(n40), .Y(n455) );
  OAI22XL U1247 ( .A0(n30), .A1(n627), .B0(n626), .B1(n28), .Y(n487) );
  CLKINVX1 U1248 ( .A(n272), .Y(n273) );
  ADDFXL U1249 ( .A(n272), .B(n440), .CI(n486), .CO(n265), .S(n266) );
  OAI22XL U1250 ( .A0(n741), .A1(n578), .B0(n46), .B1(n577), .Y(n440) );
  ADDFXL U1251 ( .A(n475), .B(n520), .CI(n305), .CO(n302), .S(n303) );
  OAI22XL U1252 ( .A0(n18), .A1(n663), .B0(n662), .B1(n16), .Y(n520) );
  OAI22XL U1253 ( .A0(n36), .A1(n615), .B0(n614), .B1(n34), .Y(n475) );
  CLKINVX1 U1254 ( .A(n304), .Y(n305) );
  ADDFXL U1255 ( .A(n304), .B(n474), .CI(n519), .CO(n294), .S(n295) );
  OAI22XL U1256 ( .A0(n36), .A1(n614), .B0(n613), .B1(n34), .Y(n474) );
  CLKINVX1 U1257 ( .A(n43), .Y(n757) );
  OAI22XL U1258 ( .A0(n742), .A1(n591), .B0(n590), .B1(n40), .Y(n252) );
  OAI22XL U1259 ( .A0(n741), .A1(n577), .B0(n46), .B1(n576), .Y(n260) );
  CMPR42X1 U1260 ( .A(n260), .B(n468), .C(n439), .D(n452), .ICI(n257), .S(n256), .ICO(n254), .CO(n255) );
  OAI22XL U1261 ( .A0(n575), .A1(n46), .B0(n741), .B1(n576), .Y(n439) );
  OAI22XL U1262 ( .A0(n592), .A1(n742), .B0(n591), .B1(n40), .Y(n452) );
  CMPR42X1 U1263 ( .A(n469), .B(n261), .C(n265), .D(n453), .ICI(n262), .S(n259), .ICO(n257), .CO(n258) );
  OAI22XL U1264 ( .A0(n36), .A1(n609), .B0(n608), .B1(n34), .Y(n469) );
  OAI22XL U1265 ( .A0(n592), .A1(n40), .B0(n593), .B1(n742), .Y(n453) );
  CLKINVX1 U1266 ( .A(n260), .Y(n261) );
  OAI22XL U1267 ( .A0(n574), .A1(n741), .B0(n46), .B1(n573), .Y(n437) );
  CLKINVX1 U1268 ( .A(n252), .Y(n253) );
  OAI22XL U1269 ( .A0(n574), .A1(n46), .B0(n575), .B1(n741), .Y(n438) );
  XNOR2X1 U1270 ( .A(n717), .B(n43), .Y(n573) );
  XNOR2X1 U1271 ( .A(b_25_), .B(n43), .Y(n572) );
  XNOR2X1 U1272 ( .A(n49), .B(n1), .Y(n714) );
  OAI22X1 U1273 ( .A0(n715), .A1(n4), .B0(n5), .B1(n764), .Y(n435) );
  CLKINVX1 U1274 ( .A(n25), .Y(n760) );
  NAND2BX1 U1275 ( .AN(n49), .B(n25), .Y(n643) );
  CMPR42X1 U1276 ( .A(n513), .B(n430), .C(n394), .D(n398), .ICI(n391), .S(n388), .ICO(n386), .CO(n387) );
  OAI22XL U1277 ( .A0(n625), .A1(n34), .B0(n36), .B1(n759), .Y(n430) );
  OAI22XL U1278 ( .A0(n656), .A1(n24), .B0(n655), .B1(n21), .Y(n513) );
  CLKINVX1 U1279 ( .A(n31), .Y(n759) );
  XNOR2X1 U1280 ( .A(n850), .B(b_15_), .Y(n686) );
  XNOR2X1 U1281 ( .A(n1), .B(b_10_), .Y(n704) );
  XNOR2X1 U1282 ( .A(n1), .B(n717), .Y(n699) );
  XNOR2X1 U1283 ( .A(n1), .B(n721), .Y(n703) );
  XNOR2X1 U1284 ( .A(n850), .B(n721), .Y(n685) );
  XNOR2X1 U1285 ( .A(n19), .B(n721), .Y(n649) );
  XNOR2X1 U1286 ( .A(n850), .B(n723), .Y(n687) );
  XNOR2X1 U1287 ( .A(n1), .B(n723), .Y(n705) );
  XNOR2X1 U1288 ( .A(n13), .B(n723), .Y(n669) );
  XNOR2X1 U1289 ( .A(n1), .B(n720), .Y(n702) );
  XNOR2X1 U1290 ( .A(n19), .B(n720), .Y(n648) );
  XNOR2X1 U1291 ( .A(n1), .B(n731), .Y(n713) );
  XNOR2X1 U1292 ( .A(n25), .B(n731), .Y(n641) );
  XNOR2X1 U1293 ( .A(n13), .B(n729), .Y(n675) );
  XNOR2X1 U1294 ( .A(n728), .B(n850), .Y(n692) );
  XNOR2X1 U1295 ( .A(n730), .B(n13), .Y(n676) );
  XNOR2X1 U1296 ( .A(n718), .B(n1), .Y(n700) );
  XNOR2X1 U1297 ( .A(b_14_), .B(n850), .Y(n689) );
  XNOR2X1 U1298 ( .A(n726), .B(n850), .Y(n690) );
  XNOR2X1 U1299 ( .A(n724), .B(n1), .Y(n706) );
  XNOR2X1 U1300 ( .A(n727), .B(n850), .Y(n691) );
  XNOR2X1 U1301 ( .A(b_7_), .B(n1), .Y(n707) );
  XNOR2X1 U1302 ( .A(n719), .B(n1), .Y(n701) );
  XNOR2X1 U1303 ( .A(n726), .B(n1), .Y(n708) );
  XNOR2X1 U1304 ( .A(n1), .B(b_16_), .Y(n698) );
  ADDHX1 U1305 ( .A(n569), .B(n434), .CO(n426), .S(n427) );
  ADDFX2 U1306 ( .A(n433), .B(n535), .CI(n423), .CO(n420), .S(n421) );
  OAI22XL U1307 ( .A0(n679), .A1(n16), .B0(n18), .B1(n762), .Y(n433) );
  OAI22XL U1308 ( .A0(n678), .A1(n17), .B0(n677), .B1(n15), .Y(n535) );
  CLKINVX1 U1309 ( .A(n13), .Y(n762) );
  CLKBUFX3 U1310 ( .A(n749), .Y(n46) );
  CLKBUFX3 U1311 ( .A(n754), .Y(n16) );
  CLKBUFX3 U1312 ( .A(n752), .Y(n28) );
  CLKBUFX3 U1313 ( .A(n750), .Y(n40) );
  CLKBUFX3 U1314 ( .A(n751), .Y(n34) );
  CLKBUFX3 U1315 ( .A(n754), .Y(n15) );
  CLKBUFX3 U1316 ( .A(n756), .Y(n4) );
  CLKBUFX3 U1317 ( .A(n746), .Y(n17) );
  CLKBUFX3 U1318 ( .A(n742), .Y(n41) );
  CLKBUFX3 U1319 ( .A(n746), .Y(n18) );
  CLKINVX1 U1320 ( .A(n19), .Y(n761) );
  CLKINVX1 U1321 ( .A(n37), .Y(n758) );
  XNOR2X1 U1322 ( .A(n19), .B(n717), .Y(n645) );
  XNOR2X1 U1323 ( .A(n19), .B(b_29_), .Y(n644) );
  NAND2X1 U1324 ( .A(n737), .B(n753), .Y(n745) );
  XOR2X1 U1325 ( .A(a_7_), .B(a_6_), .Y(n737) );
  NAND2X1 U1326 ( .A(n736), .B(n752), .Y(n744) );
  XOR2X1 U1327 ( .A(a_9_), .B(a_8_), .Y(n736) );
  NAND2X1 U1328 ( .A(n735), .B(n751), .Y(n743) );
  XOR2X1 U1329 ( .A(a_11_), .B(a_10_), .Y(n735) );
  XOR2X1 U1330 ( .A(a_13_), .B(a_12_), .Y(n734) );
  NAND2X1 U1331 ( .A(n739), .B(n755), .Y(n747) );
  XOR2X1 U1332 ( .A(a_3_), .B(a_2_), .Y(n739) );
  XOR2X1 U1333 ( .A(a_14_), .B(a_15_), .Y(n733) );
  NAND2X1 U1334 ( .A(n740), .B(n756), .Y(n748) );
  XOR2X1 U1335 ( .A(a_0_), .B(a_1_), .Y(n740) );
endmodule


module FFT_ultrafast2_shift_DW_mult_uns_9 ( a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_, 
        b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, product_31_, product_30_, 
        product_29_, product_28_, product_27_, product_26_, product_25_, 
        product_24_, product_23_, product_22_, product_21_, product_20_, 
        product_19_, product_18_, product_17_, product_16_, product_15_, 
        product_14_, product_13_, product_12_, product_11_, product_10_, 
        product_9_, product_8_, product_7_, product_6_, product_5_, product_4_, 
        product_3_, product_2_, product_1_, product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_, b_16_, b_15_, b_14_, b_13_, b_12_,
         b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_,
         b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n3, n6, n7, n9, n10, n12, n13, n15, n16, n18, n19, n21, n22, n24,
         n25, n28, n29, n31, n33, n34, n36, n37, n40, n42, n43, n45, n46, n47,
         n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n83, n84, n85, n86, n87, n89, n91, n92, n93,
         n94, n95, n97, n99, n100, n101, n102, n103, n105, n107, n108, n109,
         n110, n111, n113, n115, n116, n117, n118, n119, n121, n123, n124,
         n125, n126, n127, n129, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n178, n180, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n201, n203, n204, n205, n206, n207, n209, n211,
         n212, n213, n214, n216, n218, n220, n222, n224, n226, n228, n229,
         n230, n231, n232, n233, n235, n236, n238, n239, n240, n241, n243,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848;

  AOI21X2 U694 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  BUFX2 U695 ( .A(n742), .Y(n42) );
  OAI22X1 U696 ( .A0(n710), .A1(n748), .B0(n709), .B1(n3), .Y(n567) );
  XNOR2X1 U697 ( .A(n728), .B(n1), .Y(n710) );
  AOI21X2 U698 ( .A0(n174), .A1(n166), .B0(n167), .Y(n165) );
  OAI21X1 U699 ( .A0(n168), .A1(n172), .B0(n169), .Y(n167) );
  XNOR2X2 U700 ( .A(n724), .B(n13), .Y(n670) );
  OAI22X2 U701 ( .A0(n708), .A1(n748), .B0(n707), .B1(n3), .Y(n565) );
  XNOR2X1 U702 ( .A(n725), .B(n1), .Y(n707) );
  XNOR2X2 U703 ( .A(a_3_), .B(a_4_), .Y(n754) );
  XNOR2X2 U704 ( .A(n80), .B(n212), .Y(product_2_) );
  OAI21X2 U705 ( .A0(n173), .A1(n171), .B0(n172), .Y(n170) );
  INVX1 U706 ( .A(n174), .Y(n173) );
  ADDFX2 U707 ( .A(n547), .B(n531), .CI(n501), .CO(n403), .S(n404) );
  OAI22X1 U708 ( .A0(n674), .A1(n746), .B0(n673), .B1(n15), .Y(n531) );
  NAND2X2 U709 ( .A(n571), .B(n435), .Y(n214) );
  OAI22X1 U710 ( .A0(n715), .A1(n3), .B0(n6), .B1(n844), .Y(n435) );
  OAI22X1 U711 ( .A0(n707), .A1(n748), .B0(n706), .B1(n3), .Y(n564) );
  OAI22X1 U712 ( .A0(n714), .A1(n6), .B0(n713), .B1(n3), .Y(n571) );
  XNOR2XL U713 ( .A(n49), .B(n1), .Y(n714) );
  OAI21X4 U714 ( .A0(n127), .A1(n125), .B0(n126), .Y(n124) );
  AOI21X4 U715 ( .A0(n132), .A1(n837), .B0(n129), .Y(n127) );
  OAI22X1 U716 ( .A0(n712), .A1(n3), .B0(n6), .B1(n713), .Y(n570) );
  XNOR2X1 U717 ( .A(n7), .B(n731), .Y(n695) );
  AOI21X2 U718 ( .A0(n835), .A1(n212), .B0(n209), .Y(n207) );
  NOR2X4 U719 ( .A(n152), .B(n149), .Y(n147) );
  NAND2X1 U720 ( .A(n845), .B(n846), .Y(n712) );
  NAND2X1 U721 ( .A(n843), .B(n844), .Y(n846) );
  NAND2X1 U722 ( .A(n570), .B(n554), .Y(n211) );
  OAI22XL U723 ( .A0(n710), .A1(n3), .B0(n748), .B1(n711), .Y(n568) );
  OAI21X1 U724 ( .A0(n207), .A1(n205), .B0(n206), .Y(n204) );
  XNOR2X2 U725 ( .A(n7), .B(n729), .Y(n693) );
  XOR2X1 U726 ( .A(n79), .B(n207), .Y(product_3_) );
  OAI22XL U727 ( .A0(n661), .A1(n22), .B0(n24), .B1(n761), .Y(n432) );
  OAI22XL U728 ( .A0(n6), .A1(n705), .B0(n704), .B1(n3), .Y(n562) );
  CMPR42X1 U729 ( .A(n431), .B(n406), .C(n410), .D(n404), .ICI(n407), .S(n402), 
        .ICO(n400), .CO(n401) );
  OAI22XL U730 ( .A0(n638), .A1(n28), .B0(n29), .B1(n639), .Y(n498) );
  OR2X1 U731 ( .A(n402), .B(n408), .Y(n834) );
  ADDFXL U732 ( .A(n377), .B(n559), .CI(n482), .CO(n374), .S(n375) );
  OAI22XL U733 ( .A0(n652), .A1(n24), .B0(n651), .B1(n22), .Y(n509) );
  OAI22XL U734 ( .A0(n18), .A1(n668), .B0(n667), .B1(n16), .Y(n525) );
  OAI22XL U735 ( .A0(n18), .A1(n667), .B0(n666), .B1(n16), .Y(n524) );
  NAND2X2 U736 ( .A(n734), .B(n750), .Y(n742) );
  CLKBUFX3 U737 ( .A(n744), .Y(n29) );
  NAND2X1 U738 ( .A(n749), .B(n733), .Y(n741) );
  NOR2X1 U739 ( .A(n157), .B(n162), .Y(n155) );
  OAI21X1 U740 ( .A0(n149), .A1(n153), .B0(n150), .Y(n148) );
  CLKINVX1 U741 ( .A(n157), .Y(n233) );
  XOR2X1 U742 ( .A(n154), .B(n68), .Y(product_14_) );
  OAI22X1 U743 ( .A0(n48), .A1(n573), .B0(n46), .B1(n572), .Y(n246) );
  OAI21X1 U744 ( .A0(n111), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X1 U745 ( .A0(n103), .A1(n101), .B0(n102), .Y(n100) );
  OAI21X1 U746 ( .A0(n119), .A1(n117), .B0(n118), .Y(n116) );
  NOR2X1 U747 ( .A(n282), .B(n289), .Y(n117) );
  OAI21XL U748 ( .A0(n87), .A1(n85), .B0(n86), .Y(n84) );
  CLKINVX1 U749 ( .A(n133), .Y(n228) );
  XNOR2X1 U750 ( .A(n731), .B(n43), .Y(n587) );
  NAND2X4 U751 ( .A(n738), .B(n754), .Y(n746) );
  OAI22X1 U752 ( .A0(n692), .A1(n747), .B0(n691), .B1(n9), .Y(n549) );
  NAND2X2 U753 ( .A(n739), .B(n755), .Y(n747) );
  OR2X1 U754 ( .A(n425), .B(n426), .Y(n833) );
  OR2X1 U755 ( .A(n570), .B(n554), .Y(n835) );
  OR2X1 U756 ( .A(n290), .B(n297), .Y(n836) );
  OR2X1 U757 ( .A(n308), .B(n316), .Y(n837) );
  OR2X1 U758 ( .A(n281), .B(n276), .Y(n838) );
  OR2X1 U759 ( .A(n268), .B(n264), .Y(n839) );
  OR2X1 U760 ( .A(n256), .B(n258), .Y(n840) );
  OR2X1 U761 ( .A(n250), .B(n249), .Y(n841) );
  BUFX4 U762 ( .A(a_1_), .Y(n1) );
  BUFX4 U763 ( .A(n745), .Y(n24) );
  CLKINVX1 U764 ( .A(n184), .Y(n238) );
  BUFX4 U765 ( .A(n748), .Y(n6) );
  BUFX4 U766 ( .A(n747), .Y(n12) );
  XNOR2X1 U767 ( .A(n728), .B(n13), .Y(n674) );
  OAI22X1 U768 ( .A0(n640), .A1(n29), .B0(n639), .B1(n28), .Y(n499) );
  NOR2X2 U769 ( .A(n350), .B(n360), .Y(n149) );
  OAI21X4 U770 ( .A0(n157), .A1(n163), .B0(n158), .Y(n156) );
  NOR2X4 U771 ( .A(n370), .B(n379), .Y(n157) );
  XNOR2X1 U772 ( .A(n730), .B(n7), .Y(n694) );
  NOR2X4 U773 ( .A(n361), .B(n369), .Y(n152) );
  CMPR42X2 U774 ( .A(n374), .B(n367), .C(n372), .D(n364), .ICI(n368), .S(n361), 
        .ICO(n359), .CO(n360) );
  XNOR2X1 U775 ( .A(n727), .B(n1), .Y(n709) );
  XNOR2X1 U776 ( .A(n724), .B(n19), .Y(n652) );
  CLKBUFX4 U777 ( .A(a_7_), .Y(n19) );
  XNOR2X4 U778 ( .A(n13), .B(n721), .Y(n667) );
  CLKBUFX4 U779 ( .A(a_5_), .Y(n13) );
  CMPR42X2 U780 ( .A(n393), .B(n499), .C(n529), .D(n484), .ICI(n397), .S(n391), 
        .ICO(n389), .CO(n390) );
  ADDHX1 U781 ( .A(n561), .B(n545), .CO(n392), .S(n393) );
  XNOR2X1 U782 ( .A(n727), .B(n13), .Y(n673) );
  NOR2BX1 U783 ( .AN(n49), .B(n9), .Y(n554) );
  CLKBUFX4 U784 ( .A(a_3_), .Y(n7) );
  XOR2X1 U785 ( .A(n199), .B(n77), .Y(product_5_) );
  ADDHX1 U786 ( .A(n563), .B(n515), .CO(n405), .S(n406) );
  OAI22X1 U787 ( .A0(n697), .A1(n10), .B0(n12), .B1(n763), .Y(n434) );
  AND2X1 U788 ( .A(n164), .B(n155), .Y(n842) );
  NOR2X4 U789 ( .A(n842), .B(n156), .Y(n154) );
  NAND2XL U790 ( .A(n730), .B(n1), .Y(n845) );
  INVXL U791 ( .A(n730), .Y(n843) );
  INVXL U792 ( .A(n1), .Y(n844) );
  BUFX8 U793 ( .A(b_2_), .Y(n730) );
  OAI22X1 U794 ( .A0(n712), .A1(n6), .B0(n711), .B1(n3), .Y(n569) );
  XOR2X1 U795 ( .A(n135), .B(n64), .Y(product_18_) );
  INVX3 U796 ( .A(n165), .Y(n164) );
  CLKBUFX2 U797 ( .A(b_8_), .Y(n724) );
  ADDFX2 U798 ( .A(n502), .B(n564), .CI(n532), .CO(n410), .S(n411) );
  XNOR2X1 U799 ( .A(n37), .B(n729), .Y(n603) );
  XNOR2XL U800 ( .A(n19), .B(n723), .Y(n651) );
  BUFX3 U801 ( .A(n743), .Y(n36) );
  OAI21X2 U802 ( .A0(n145), .A1(n165), .B0(n146), .Y(n144) );
  CLKBUFX2 U803 ( .A(b_7_), .Y(n725) );
  OAI21X1 U804 ( .A0(n154), .A1(n152), .B0(n153), .Y(n151) );
  CLKBUFX2 U805 ( .A(b_5_), .Y(n727) );
  OAI22X1 U806 ( .A0(n676), .A1(n746), .B0(n675), .B1(n15), .Y(n533) );
  CLKINVX1 U807 ( .A(n131), .Y(n129) );
  AOI21X1 U808 ( .A0(n92), .A1(n841), .B0(n89), .Y(n87) );
  NOR2X1 U809 ( .A(n190), .B(n193), .Y(n188) );
  XNOR2XL U810 ( .A(n725), .B(n19), .Y(n653) );
  XNOR2XL U811 ( .A(n726), .B(n19), .Y(n654) );
  XNOR2XL U812 ( .A(n37), .B(n731), .Y(n605) );
  XNOR2XL U813 ( .A(n31), .B(n729), .Y(n621) );
  INVX1 U814 ( .A(a_0_), .Y(n756) );
  NAND2XL U815 ( .A(n232), .B(n153), .Y(n68) );
  INVXL U816 ( .A(n149), .Y(n231) );
  XNOR2X1 U817 ( .A(n19), .B(n729), .Y(n657) );
  XNOR2X1 U818 ( .A(n724), .B(n7), .Y(n688) );
  NOR2XL U819 ( .A(n141), .B(n138), .Y(n136) );
  OAI21X1 U820 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NAND2X1 U821 ( .A(n425), .B(n426), .Y(n203) );
  NOR2BXL U822 ( .AN(n49), .B(n33), .Y(n485) );
  XNOR2XL U823 ( .A(n13), .B(n731), .Y(n677) );
  XNOR2XL U824 ( .A(n19), .B(n731), .Y(n659) );
  XNOR2XL U825 ( .A(n13), .B(n722), .Y(n668) );
  INVXL U826 ( .A(n138), .Y(n229) );
  OAI21XL U827 ( .A0(n138), .A1(n142), .B0(n139), .Y(n137) );
  NAND2XL U828 ( .A(n836), .B(n123), .Y(n61) );
  NAND2X1 U829 ( .A(n238), .B(n185), .Y(n74) );
  CLKINVX1 U830 ( .A(n185), .Y(n183) );
  XOR2X1 U831 ( .A(n173), .B(n72), .Y(product_10_) );
  INVXL U832 ( .A(n193), .Y(n240) );
  OAI22X1 U833 ( .A0(n642), .A1(n29), .B0(n641), .B1(n28), .Y(n501) );
  OAI22XL U834 ( .A0(n622), .A1(n36), .B0(n621), .B1(n33), .Y(n482) );
  XNOR2X1 U835 ( .A(n730), .B(n19), .Y(n658) );
  XNOR2X1 U836 ( .A(n49), .B(n19), .Y(n660) );
  CLKBUFX3 U837 ( .A(a_15_), .Y(n43) );
  INVXL U838 ( .A(n7), .Y(n763) );
  OAI21X1 U839 ( .A0(n143), .A1(n141), .B0(n142), .Y(n140) );
  CLKBUFX2 U840 ( .A(b_14_), .Y(n718) );
  CLKBUFX4 U841 ( .A(b_0_), .Y(n49) );
  NAND2XL U842 ( .A(n233), .B(n158), .Y(n69) );
  OAI21X2 U843 ( .A0(n95), .A1(n93), .B0(n94), .Y(n92) );
  NAND2XL U844 ( .A(n835), .B(n211), .Y(n80) );
  CLKBUFX2 U845 ( .A(b_6_), .Y(n726) );
  CLKBUFX2 U846 ( .A(b_1_), .Y(n731) );
  INVXL U847 ( .A(n187), .Y(n186) );
  NOR2X1 U848 ( .A(n339), .B(n349), .Y(n141) );
  NOR2X1 U849 ( .A(n328), .B(n338), .Y(n138) );
  NOR2X1 U850 ( .A(n317), .B(n327), .Y(n133) );
  NOR2X1 U851 ( .A(n298), .B(n307), .Y(n125) );
  OAI21X2 U852 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  NAND2XL U853 ( .A(n235), .B(n169), .Y(n71) );
  INVXL U854 ( .A(n168), .Y(n235) );
  NOR2X1 U855 ( .A(n409), .B(n413), .Y(n184) );
  NAND2XL U856 ( .A(n243), .B(n206), .Y(n79) );
  NAND2XL U857 ( .A(n241), .B(n198), .Y(n77) );
  NAND2XL U858 ( .A(n236), .B(n172), .Y(n72) );
  NAND2XL U859 ( .A(n240), .B(n194), .Y(n76) );
  XNOR2XL U860 ( .A(n164), .B(n70), .Y(product_12_) );
  NAND2XL U861 ( .A(n160), .B(n163), .Y(n70) );
  INVXL U862 ( .A(n190), .Y(n239) );
  XNOR2XL U863 ( .A(n204), .B(n78), .Y(product_4_) );
  XNOR2X1 U864 ( .A(n847), .B(n73), .Y(product_9_) );
  AO21XL U865 ( .A0(n186), .A1(n238), .B0(n183), .Y(n847) );
  NAND2XL U866 ( .A(n414), .B(n418), .Y(n191) );
  INVXL U867 ( .A(n163), .Y(n161) );
  NOR2X1 U868 ( .A(n275), .B(n269), .Y(n109) );
  NOR2X1 U869 ( .A(n263), .B(n259), .Y(n101) );
  NOR2X1 U870 ( .A(n255), .B(n251), .Y(n93) );
  NOR2X1 U871 ( .A(n248), .B(n247), .Y(n85) );
  ADDHX1 U872 ( .A(n533), .B(n549), .CO(n415), .S(n416) );
  NOR2BXL U873 ( .AN(n49), .B(n28), .Y(n502) );
  OAI22X1 U874 ( .A0(n690), .A1(n12), .B0(n689), .B1(n9), .Y(n547) );
  NOR2BXL U875 ( .AN(n49), .B(n15), .Y(n536) );
  CMPR42X2 U876 ( .A(n497), .B(n381), .C(n382), .D(n373), .ICI(n378), .S(n370), 
        .ICO(n368), .CO(n369) );
  NOR2X1 U877 ( .A(n380), .B(n387), .Y(n162) );
  XNOR2XL U878 ( .A(n49), .B(n43), .Y(n588) );
  NOR2X1 U879 ( .A(n396), .B(n401), .Y(n171) );
  NOR2X1 U880 ( .A(n419), .B(n420), .Y(n193) );
  NOR2BXL U881 ( .AN(n49), .B(n45), .Y(n450) );
  NOR2X1 U882 ( .A(n427), .B(n553), .Y(n205) );
  NOR2X1 U883 ( .A(n421), .B(n424), .Y(n197) );
  NAND2BXL U884 ( .AN(n213), .B(n214), .Y(n81) );
  NOR2XL U885 ( .A(n571), .B(n435), .Y(n213) );
  XNOR2XL U886 ( .A(n730), .B(n43), .Y(n586) );
  NOR2BXL U887 ( .AN(n49), .B(n3), .Y(product_0_) );
  NAND2BXL U888 ( .AN(n49), .B(n43), .Y(n589) );
  XNOR2XL U889 ( .A(n727), .B(n43), .Y(n583) );
  XNOR2XL U890 ( .A(n726), .B(n43), .Y(n582) );
  XNOR2XL U891 ( .A(n725), .B(n43), .Y(n581) );
  XNOR2XL U892 ( .A(n724), .B(n43), .Y(n580) );
  XNOR2XL U893 ( .A(n728), .B(n43), .Y(n584) );
  XNOR2XL U894 ( .A(n729), .B(n43), .Y(n585) );
  OAI22XL U895 ( .A0(n24), .A1(n649), .B0(n648), .B1(n22), .Y(n324) );
  OAI22XL U896 ( .A0(n24), .A1(n645), .B0(n644), .B1(n22), .Y(n286) );
  AO21XL U897 ( .A0(n18), .A1(n16), .B0(n662), .Y(n519) );
  AO21XL U898 ( .A0(n6), .A1(n756), .B0(n698), .Y(n555) );
  AO21XL U899 ( .A0(n12), .A1(n10), .B0(n680), .Y(n537) );
  AO21XL U900 ( .A0(n24), .A1(n22), .B0(n644), .Y(n503) );
  XNOR2XL U901 ( .A(n719), .B(n43), .Y(n575) );
  XNOR2XL U902 ( .A(n718), .B(n43), .Y(n574) );
  XNOR2XL U903 ( .A(n723), .B(n43), .Y(n579) );
  XNOR2XL U904 ( .A(n722), .B(n43), .Y(n578) );
  XNOR2XL U905 ( .A(n721), .B(n43), .Y(n577) );
  XNOR2XL U906 ( .A(n43), .B(n720), .Y(n576) );
  AO21XL U907 ( .A0(n744), .A1(n28), .B0(n626), .Y(n486) );
  AO21XL U908 ( .A0(n36), .A1(n34), .B0(n608), .Y(n468) );
  ADDFXL U909 ( .A(n253), .B(n438), .CI(n254), .CO(n250), .S(n251) );
  ADDFXL U910 ( .A(n252), .B(n451), .CI(n437), .CO(n248), .S(n249) );
  AO21XL U911 ( .A0(n42), .A1(n40), .B0(n590), .Y(n451) );
  AO21XL U912 ( .A0(n48), .A1(n46), .B0(n572), .Y(n436) );
  XNOR2XL U913 ( .A(n49), .B(n7), .Y(n696) );
  NAND2BXL U914 ( .AN(n49), .B(n1), .Y(n715) );
  XNOR2XL U915 ( .A(n725), .B(n13), .Y(n671) );
  XNOR2XL U916 ( .A(n725), .B(n25), .Y(n635) );
  XNOR2XL U917 ( .A(n719), .B(n7), .Y(n683) );
  XNOR2XL U918 ( .A(n726), .B(n13), .Y(n672) );
  XNOR2XL U919 ( .A(n726), .B(n25), .Y(n636) );
  XNOR2XL U920 ( .A(n727), .B(n25), .Y(n637) );
  XNOR2XL U921 ( .A(n727), .B(n31), .Y(n619) );
  XNOR2XL U922 ( .A(n727), .B(n19), .Y(n655) );
  XNOR2XL U923 ( .A(n728), .B(n25), .Y(n638) );
  XNOR2XL U924 ( .A(n728), .B(n19), .Y(n656) );
  XNOR2XL U925 ( .A(n728), .B(n31), .Y(n620) );
  XNOR2XL U926 ( .A(n730), .B(n25), .Y(n640) );
  XNOR2XL U927 ( .A(n730), .B(n31), .Y(n622) );
  XNOR2XL U928 ( .A(n730), .B(n37), .Y(n604) );
  XNOR2XL U929 ( .A(n31), .B(n731), .Y(n623) );
  XNOR2XL U930 ( .A(n1), .B(n729), .Y(n711) );
  XNOR2XL U931 ( .A(n49), .B(n25), .Y(n642) );
  XNOR2XL U932 ( .A(n49), .B(n13), .Y(n678) );
  XNOR2XL U933 ( .A(n49), .B(n31), .Y(n624) );
  XNOR2XL U934 ( .A(n49), .B(n37), .Y(n606) );
  NAND2BXL U935 ( .AN(n49), .B(n7), .Y(n697) );
  NAND2BXL U936 ( .AN(n49), .B(n19), .Y(n661) );
  NAND2BXL U937 ( .AN(n49), .B(n13), .Y(n679) );
  NAND2BXL U938 ( .AN(n49), .B(n37), .Y(n607) );
  XNOR2XL U939 ( .A(n725), .B(n31), .Y(n617) );
  XNOR2XL U940 ( .A(n724), .B(n25), .Y(n634) );
  XNOR2XL U941 ( .A(n719), .B(n13), .Y(n665) );
  XNOR2XL U942 ( .A(n726), .B(n31), .Y(n618) );
  XNOR2XL U943 ( .A(n727), .B(n37), .Y(n601) );
  XNOR2XL U944 ( .A(n724), .B(n31), .Y(n616) );
  XNOR2XL U945 ( .A(n726), .B(n37), .Y(n600) );
  XNOR2XL U946 ( .A(n718), .B(n7), .Y(n682) );
  XNOR2XL U947 ( .A(n728), .B(n37), .Y(n602) );
  XNOR2XL U948 ( .A(n718), .B(n13), .Y(n664) );
  XNOR2XL U949 ( .A(n19), .B(n722), .Y(n650) );
  XNOR2XL U950 ( .A(n25), .B(n729), .Y(n639) );
  XNOR2XL U951 ( .A(n7), .B(n720), .Y(n684) );
  XNOR2XL U952 ( .A(n13), .B(n720), .Y(n666) );
  NAND2BXL U953 ( .AN(n49), .B(n31), .Y(n625) );
  XNOR2XL U954 ( .A(n719), .B(n19), .Y(n647) );
  XNOR2XL U955 ( .A(n725), .B(n37), .Y(n599) );
  XNOR2XL U956 ( .A(n724), .B(n37), .Y(n598) );
  XNOR2XL U957 ( .A(n719), .B(n25), .Y(n629) );
  XNOR2XL U958 ( .A(n719), .B(n31), .Y(n611) );
  XNOR2XL U959 ( .A(n718), .B(n19), .Y(n646) );
  XNOR2XL U960 ( .A(n718), .B(n25), .Y(n628) );
  XNOR2XL U961 ( .A(n718), .B(n31), .Y(n610) );
  XNOR2XL U962 ( .A(n7), .B(n717), .Y(n681) );
  XNOR2XL U963 ( .A(n25), .B(n722), .Y(n632) );
  XNOR2XL U964 ( .A(n13), .B(n717), .Y(n663) );
  XNOR2XL U965 ( .A(n31), .B(n722), .Y(n614) );
  XNOR2XL U966 ( .A(n37), .B(n722), .Y(n596) );
  XNOR2XL U967 ( .A(n25), .B(n723), .Y(n633) );
  XNOR2XL U968 ( .A(n31), .B(n723), .Y(n615) );
  XNOR2XL U969 ( .A(n37), .B(n723), .Y(n597) );
  XNOR2XL U970 ( .A(n25), .B(n721), .Y(n631) );
  XNOR2XL U971 ( .A(n31), .B(n721), .Y(n613) );
  XNOR2XL U972 ( .A(n37), .B(n721), .Y(n595) );
  XNOR2XL U973 ( .A(n25), .B(n720), .Y(n630) );
  XNOR2XL U974 ( .A(n31), .B(n720), .Y(n612) );
  XNOR2XL U975 ( .A(n7), .B(n716), .Y(n680) );
  XNOR2XL U976 ( .A(n13), .B(n716), .Y(n662) );
  XNOR2XL U977 ( .A(n719), .B(n37), .Y(n593) );
  XNOR2XL U978 ( .A(n718), .B(n37), .Y(n592) );
  XNOR2XL U979 ( .A(n25), .B(n717), .Y(n627) );
  XNOR2XL U980 ( .A(n37), .B(n720), .Y(n594) );
  XNOR2XL U981 ( .A(n25), .B(n716), .Y(n626) );
  XNOR2XL U982 ( .A(n31), .B(n717), .Y(n609) );
  XNOR2XL U983 ( .A(n37), .B(n717), .Y(n591) );
  XNOR2XL U984 ( .A(n31), .B(n716), .Y(n608) );
  XNOR2XL U985 ( .A(n37), .B(n716), .Y(n590) );
  XNOR2X1 U986 ( .A(a_5_), .B(a_6_), .Y(n753) );
  XNOR2X1 U987 ( .A(a_1_), .B(a_2_), .Y(n755) );
  XNOR2X1 U988 ( .A(a_7_), .B(a_8_), .Y(n752) );
  XNOR2X1 U989 ( .A(a_11_), .B(a_12_), .Y(n750) );
  XNOR2X1 U990 ( .A(a_9_), .B(a_10_), .Y(n751) );
  CLKBUFX3 U991 ( .A(a_9_), .Y(n25) );
  CLKBUFX3 U992 ( .A(a_11_), .Y(n31) );
  CLKBUFX3 U993 ( .A(a_13_), .Y(n37) );
  XNOR2X1 U994 ( .A(a_13_), .B(a_14_), .Y(n749) );
  XNOR2X1 U995 ( .A(n140), .B(n65), .Y(product_17_) );
  NAND2X1 U996 ( .A(n229), .B(n139), .Y(n65) );
  XNOR2X1 U997 ( .A(n132), .B(n63), .Y(product_19_) );
  NAND2X1 U998 ( .A(n837), .B(n131), .Y(n63) );
  AOI21X1 U999 ( .A0(n144), .A1(n136), .B0(n137), .Y(n135) );
  OAI21X1 U1000 ( .A0(n135), .A1(n133), .B0(n134), .Y(n132) );
  XOR2X1 U1001 ( .A(n127), .B(n62), .Y(product_20_) );
  NAND2X1 U1002 ( .A(n226), .B(n126), .Y(n62) );
  CLKINVX1 U1003 ( .A(n125), .Y(n226) );
  NAND2X1 U1004 ( .A(n228), .B(n134), .Y(n64) );
  XOR2X1 U1005 ( .A(n143), .B(n66), .Y(product_16_) );
  NAND2X1 U1006 ( .A(n230), .B(n142), .Y(n66) );
  CLKINVX1 U1007 ( .A(n141), .Y(n230) );
  CLKINVX1 U1008 ( .A(n144), .Y(n143) );
  XNOR2X1 U1009 ( .A(n186), .B(n74), .Y(product_8_) );
  XNOR2X1 U1010 ( .A(n151), .B(n67), .Y(product_15_) );
  NAND2X1 U1011 ( .A(n231), .B(n150), .Y(n67) );
  XNOR2X1 U1012 ( .A(n92), .B(n53), .Y(product_29_) );
  NAND2X1 U1013 ( .A(n841), .B(n91), .Y(n53) );
  XNOR2X1 U1014 ( .A(n100), .B(n55), .Y(product_27_) );
  NAND2X1 U1015 ( .A(n840), .B(n99), .Y(n55) );
  XNOR2X1 U1016 ( .A(n108), .B(n57), .Y(product_25_) );
  NAND2X1 U1017 ( .A(n839), .B(n107), .Y(n57) );
  XNOR2X1 U1018 ( .A(n116), .B(n59), .Y(product_23_) );
  NAND2X1 U1019 ( .A(n838), .B(n115), .Y(n59) );
  XNOR2X1 U1020 ( .A(n124), .B(n61), .Y(product_21_) );
  NAND2X1 U1021 ( .A(n147), .B(n155), .Y(n145) );
  AOI21X1 U1022 ( .A0(n156), .A1(n147), .B0(n148), .Y(n146) );
  AOI21X1 U1023 ( .A0(n124), .A1(n836), .B0(n121), .Y(n119) );
  CLKINVX1 U1024 ( .A(n123), .Y(n121) );
  AOI21X1 U1025 ( .A0(n116), .A1(n838), .B0(n113), .Y(n111) );
  CLKINVX1 U1026 ( .A(n115), .Y(n113) );
  AOI21X1 U1027 ( .A0(n108), .A1(n839), .B0(n105), .Y(n103) );
  CLKINVX1 U1028 ( .A(n107), .Y(n105) );
  AOI21X1 U1029 ( .A0(n100), .A1(n840), .B0(n97), .Y(n95) );
  CLKINVX1 U1030 ( .A(n99), .Y(n97) );
  CLKINVX1 U1031 ( .A(n91), .Y(n89) );
  CLKINVX1 U1032 ( .A(n211), .Y(n209) );
  CLKBUFX3 U1033 ( .A(b_10_), .Y(n722) );
  CLKBUFX3 U1034 ( .A(b_15_), .Y(n717) );
  CLKBUFX3 U1035 ( .A(b_11_), .Y(n721) );
  CLKBUFX3 U1036 ( .A(b_4_), .Y(n728) );
  CLKBUFX3 U1037 ( .A(b_13_), .Y(n719) );
  NAND2X1 U1038 ( .A(n339), .B(n349), .Y(n142) );
  NAND2X1 U1039 ( .A(n308), .B(n316), .Y(n131) );
  NAND2X1 U1040 ( .A(n350), .B(n360), .Y(n150) );
  NAND2X1 U1041 ( .A(n328), .B(n338), .Y(n139) );
  NAND2X1 U1042 ( .A(n317), .B(n327), .Y(n134) );
  XOR2X1 U1043 ( .A(n159), .B(n69), .Y(product_13_) );
  AOI21X1 U1044 ( .A0(n164), .A1(n160), .B0(n161), .Y(n159) );
  CLKINVX1 U1045 ( .A(n152), .Y(n232) );
  XOR2X1 U1046 ( .A(n87), .B(n52), .Y(product_30_) );
  NAND2X1 U1047 ( .A(n216), .B(n86), .Y(n52) );
  CLKINVX1 U1048 ( .A(n85), .Y(n216) );
  XOR2X1 U1049 ( .A(n95), .B(n54), .Y(product_28_) );
  NAND2X1 U1050 ( .A(n218), .B(n94), .Y(n54) );
  CLKINVX1 U1051 ( .A(n93), .Y(n218) );
  XOR2X1 U1052 ( .A(n103), .B(n56), .Y(product_26_) );
  NAND2X1 U1053 ( .A(n220), .B(n102), .Y(n56) );
  CLKINVX1 U1054 ( .A(n101), .Y(n220) );
  XOR2X1 U1055 ( .A(n111), .B(n58), .Y(product_24_) );
  NAND2X1 U1056 ( .A(n222), .B(n110), .Y(n58) );
  CLKINVX1 U1057 ( .A(n109), .Y(n222) );
  XOR2X1 U1058 ( .A(n119), .B(n60), .Y(product_22_) );
  NAND2X1 U1059 ( .A(n224), .B(n118), .Y(n60) );
  CLKINVX1 U1060 ( .A(n117), .Y(n224) );
  CLKINVX1 U1061 ( .A(n196), .Y(n195) );
  NAND2X1 U1062 ( .A(n298), .B(n307), .Y(n126) );
  NAND2X1 U1063 ( .A(n833), .B(n203), .Y(n78) );
  XNOR2X1 U1064 ( .A(n170), .B(n71), .Y(product_11_) );
  XNOR2X1 U1065 ( .A(n84), .B(n51), .Y(product_31_) );
  NAND2X1 U1066 ( .A(n848), .B(n83), .Y(n51) );
  NAND2X1 U1067 ( .A(n436), .B(n246), .Y(n83) );
  CMPR42X1 U1068 ( .A(n344), .B(n334), .C(n341), .D(n331), .ICI(n337), .S(n328), .ICO(n326), .CO(n327) );
  CMPR42X1 U1069 ( .A(n366), .B(n356), .C(n363), .D(n353), .ICI(n359), .S(n350), .ICO(n348), .CO(n349) );
  CMPR42X1 U1070 ( .A(n345), .B(n355), .C(n352), .D(n342), .ICI(n348), .S(n339), .ICO(n337), .CO(n338) );
  CMPR42X1 U1071 ( .A(n318), .B(n314), .C(n311), .D(n319), .ICI(n315), .S(n308), .ICO(n306), .CO(n307) );
  CMPR42X1 U1072 ( .A(n329), .B(n333), .C(n330), .D(n320), .ICI(n326), .S(n317), .ICO(n315), .CO(n316) );
  CMPR42X1 U1073 ( .A(n303), .B(n309), .C(n310), .D(n301), .ICI(n306), .S(n298), .ICO(n296), .CO(n297) );
  OAI21X1 U1074 ( .A0(n187), .A1(n175), .B0(n176), .Y(n174) );
  NAND2X1 U1075 ( .A(n834), .B(n238), .Y(n175) );
  AOI21X1 U1076 ( .A0(n834), .A1(n183), .B0(n178), .Y(n176) );
  NOR2X1 U1077 ( .A(n168), .B(n171), .Y(n166) );
  NOR2X1 U1078 ( .A(n414), .B(n418), .Y(n190) );
  AOI21X1 U1079 ( .A0(n204), .A1(n833), .B0(n201), .Y(n199) );
  CLKINVX1 U1080 ( .A(n203), .Y(n201) );
  XNOR2X1 U1081 ( .A(n192), .B(n75), .Y(product_7_) );
  NAND2X1 U1082 ( .A(n239), .B(n191), .Y(n75) );
  OAI21XL U1083 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2X1 U1084 ( .A(n361), .B(n369), .Y(n153) );
  NAND2X1 U1085 ( .A(n409), .B(n413), .Y(n185) );
  NAND2X1 U1086 ( .A(n370), .B(n379), .Y(n158) );
  NAND2X1 U1087 ( .A(n834), .B(n180), .Y(n73) );
  CLKINVX1 U1088 ( .A(n197), .Y(n241) );
  CLKINVX1 U1089 ( .A(n205), .Y(n243) );
  XOR2X1 U1090 ( .A(n195), .B(n76), .Y(product_6_) );
  CLKINVX1 U1091 ( .A(n171), .Y(n236) );
  CLKINVX1 U1092 ( .A(n214), .Y(n212) );
  CLKINVX1 U1093 ( .A(n324), .Y(n325) );
  CLKINVX1 U1094 ( .A(n162), .Y(n160) );
  CLKINVX1 U1095 ( .A(n180), .Y(n178) );
  NAND2X1 U1096 ( .A(n281), .B(n276), .Y(n115) );
  NAND2X1 U1097 ( .A(n268), .B(n264), .Y(n107) );
  NAND2X1 U1098 ( .A(n290), .B(n297), .Y(n123) );
  NAND2X1 U1099 ( .A(n275), .B(n269), .Y(n110) );
  NAND2X1 U1100 ( .A(n282), .B(n289), .Y(n118) );
  CLKINVX1 U1101 ( .A(n286), .Y(n287) );
  NAND2X1 U1102 ( .A(n256), .B(n258), .Y(n99) );
  NAND2X1 U1103 ( .A(n263), .B(n259), .Y(n102) );
  NAND2X1 U1104 ( .A(n250), .B(n249), .Y(n91) );
  NAND2X1 U1105 ( .A(n255), .B(n251), .Y(n94) );
  NAND2X1 U1106 ( .A(n248), .B(n247), .Y(n86) );
  CLKINVX1 U1107 ( .A(n246), .Y(n247) );
  OR2X1 U1108 ( .A(n436), .B(n246), .Y(n848) );
  CMPR42X1 U1109 ( .A(n518), .B(n550), .C(n534), .D(n566), .ICI(n422), .S(n419), .ICO(n417), .CO(n418) );
  OAI22XL U1110 ( .A0(n709), .A1(n6), .B0(n708), .B1(n3), .Y(n566) );
  OAI22XL U1111 ( .A0(n676), .A1(n15), .B0(n746), .B1(n677), .Y(n534) );
  NOR2BX1 U1112 ( .AN(n49), .B(n21), .Y(n518) );
  CMPR42X1 U1113 ( .A(n516), .B(n548), .C(n415), .D(n411), .ICI(n412), .S(n409), .ICO(n407), .CO(n408) );
  OAI22XL U1114 ( .A0(n691), .A1(n747), .B0(n690), .B1(n9), .Y(n548) );
  OAI22XL U1115 ( .A0(n658), .A1(n21), .B0(n24), .B1(n659), .Y(n516) );
  CMPR42X1 U1116 ( .A(n565), .B(n432), .C(n517), .D(n416), .ICI(n417), .S(n414), .ICO(n412), .CO(n413) );
  OAI22XL U1117 ( .A0(n660), .A1(n24), .B0(n659), .B1(n21), .Y(n517) );
  OAI22XL U1118 ( .A0(n638), .A1(n29), .B0(n637), .B1(n752), .Y(n497) );
  CMPR42X1 U1119 ( .A(n528), .B(n385), .C(n390), .D(n383), .ICI(n386), .S(n380), .ICO(n378), .CO(n379) );
  OAI22XL U1120 ( .A0(n671), .A1(n746), .B0(n670), .B1(n15), .Y(n528) );
  OAI22XL U1121 ( .A0(n24), .A1(n650), .B0(n649), .B1(n22), .Y(n507) );
  NOR2X2 U1122 ( .A(n388), .B(n395), .Y(n168) );
  CLKBUFX3 U1123 ( .A(b_12_), .Y(n720) );
  CLKBUFX3 U1124 ( .A(b_3_), .Y(n729) );
  CLKBUFX3 U1125 ( .A(b_9_), .Y(n723) );
  CLKBUFX3 U1126 ( .A(b_16_), .Y(n716) );
  OAI22XL U1127 ( .A0(n692), .A1(n9), .B0(n747), .B1(n693), .Y(n550) );
  OAI22XL U1128 ( .A0(n700), .A1(n6), .B0(n699), .B1(n3), .Y(n557) );
  OAI22XL U1129 ( .A0(n682), .A1(n12), .B0(n681), .B1(n10), .Y(n539) );
  OAI22XL U1130 ( .A0(n700), .A1(n3), .B0(n701), .B1(n6), .Y(n558) );
  OAI22XL U1131 ( .A0(n29), .A1(n633), .B0(n632), .B1(n28), .Y(n492) );
  OAI22XL U1132 ( .A0(n689), .A1(n12), .B0(n688), .B1(n9), .Y(n546) );
  ADDFX2 U1133 ( .A(n536), .B(n568), .CI(n552), .CO(n424), .S(n425) );
  OAI22XL U1134 ( .A0(n694), .A1(n9), .B0(n747), .B1(n695), .Y(n552) );
  OAI22XL U1135 ( .A0(n706), .A1(n748), .B0(n705), .B1(n3), .Y(n563) );
  OAI22XL U1136 ( .A0(n658), .A1(n24), .B0(n657), .B1(n21), .Y(n515) );
  ADDHXL U1137 ( .A(n524), .B(n556), .CO(n346), .S(n347) );
  OAI22XL U1138 ( .A0(n6), .A1(n699), .B0(n698), .B1(n3), .Y(n556) );
  OAI22XL U1139 ( .A0(n6), .A1(n704), .B0(n703), .B1(n3), .Y(n561) );
  OAI22XL U1140 ( .A0(n688), .A1(n12), .B0(n687), .B1(n10), .Y(n545) );
  ADDHXL U1141 ( .A(n525), .B(n509), .CO(n357), .S(n358) );
  NAND2X1 U1142 ( .A(n380), .B(n387), .Y(n163) );
  NAND2X1 U1143 ( .A(n396), .B(n401), .Y(n172) );
  CMPR42X1 U1144 ( .A(n358), .B(n541), .C(n464), .D(n449), .ICI(n362), .S(n356), .ICO(n354), .CO(n355) );
  OAI22XL U1145 ( .A0(n683), .A1(n10), .B0(n12), .B1(n684), .Y(n541) );
  OAI22XL U1146 ( .A0(n588), .A1(n47), .B0(n45), .B1(n587), .Y(n449) );
  OAI22XL U1147 ( .A0(n604), .A1(n42), .B0(n603), .B1(n40), .Y(n464) );
  CMPR42X1 U1148 ( .A(n491), .B(n324), .C(n537), .D(n476), .ICI(n445), .S(n314), .ICO(n312), .CO(n313) );
  OAI22XL U1149 ( .A0(n616), .A1(n743), .B0(n615), .B1(n34), .Y(n476) );
  OAI22XL U1150 ( .A0(n584), .A1(n47), .B0(n583), .B1(n45), .Y(n445) );
  CMPR42X1 U1151 ( .A(n493), .B(n346), .C(n523), .D(n336), .ICI(n343), .S(n334), .ICO(n332), .CO(n333) );
  OAI22XL U1152 ( .A0(n634), .A1(n29), .B0(n633), .B1(n28), .Y(n493) );
  XNOR2X1 U1153 ( .A(n555), .B(n507), .Y(n336) );
  OAI22XL U1154 ( .A0(n665), .A1(n16), .B0(n18), .B1(n666), .Y(n523) );
  CMPR42X1 U1155 ( .A(n542), .B(n526), .C(n376), .D(n450), .ICI(n496), .S(n367), .ICO(n365), .CO(n366) );
  OAI22XL U1156 ( .A0(n637), .A1(n29), .B0(n636), .B1(n28), .Y(n496) );
  OAI22XL U1157 ( .A0(n18), .A1(n669), .B0(n668), .B1(n16), .Y(n526) );
  OAI22XL U1158 ( .A0(n12), .A1(n685), .B0(n684), .B1(n10), .Y(n542) );
  NAND2X1 U1159 ( .A(n419), .B(n420), .Y(n194) );
  CMPR42X1 U1160 ( .A(n508), .B(n347), .C(n357), .D(n540), .ICI(n479), .S(n345), .ICO(n343), .CO(n344) );
  OAI22XL U1161 ( .A0(n619), .A1(n743), .B0(n618), .B1(n33), .Y(n479) );
  OAI22XL U1162 ( .A0(n24), .A1(n651), .B0(n650), .B1(n22), .Y(n508) );
  OAI22XL U1163 ( .A0(n682), .A1(n10), .B0(n683), .B1(n12), .Y(n540) );
  NAND2X1 U1164 ( .A(n402), .B(n408), .Y(n180) );
  CMPR42X1 U1165 ( .A(n506), .B(n321), .C(n521), .D(n460), .ICI(n322), .S(n311), .ICO(n309), .CO(n310) );
  OAI22XL U1166 ( .A0(n600), .A1(n742), .B0(n599), .B1(n40), .Y(n460) );
  OAI22XL U1167 ( .A0(n664), .A1(n18), .B0(n663), .B1(n16), .Y(n521) );
  OAI22XL U1168 ( .A0(n647), .A1(n22), .B0(n24), .B1(n648), .Y(n506) );
  CMPR42X1 U1169 ( .A(n500), .B(n405), .C(n403), .D(n400), .ICI(n399), .S(n396), .ICO(n394), .CO(n395) );
  OAI22XL U1170 ( .A0(n640), .A1(n28), .B0(n29), .B1(n641), .Y(n500) );
  OAI22XL U1171 ( .A0(n624), .A1(n36), .B0(n623), .B1(n33), .Y(n484) );
  OAI22XL U1172 ( .A0(n672), .A1(n746), .B0(n671), .B1(n15), .Y(n529) );
  CMPR42X1 U1173 ( .A(n467), .B(n498), .C(n483), .D(n512), .ICI(n389), .S(n383), .ICO(n381), .CO(n382) );
  OAI22XL U1174 ( .A0(n655), .A1(n24), .B0(n654), .B1(n21), .Y(n512) );
  OAI22XL U1175 ( .A0(n622), .A1(n33), .B0(n36), .B1(n623), .Y(n483) );
  NOR2BX1 U1176 ( .AN(n49), .B(n40), .Y(n467) );
  CMPR42X1 U1177 ( .A(n494), .B(n463), .C(n448), .D(n354), .ICI(n351), .S(n342), .ICO(n340), .CO(n341) );
  OAI22XL U1178 ( .A0(n586), .A1(n45), .B0(n47), .B1(n587), .Y(n448) );
  OAI22XL U1179 ( .A0(n602), .A1(n40), .B0(n742), .B1(n603), .Y(n463) );
  OAI22XL U1180 ( .A0(n635), .A1(n29), .B0(n634), .B1(n28), .Y(n494) );
  CMPR42X1 U1181 ( .A(n558), .B(n510), .C(n481), .D(n465), .ICI(n371), .S(n364), .ICO(n362), .CO(n363) );
  OAI22XL U1182 ( .A0(n604), .A1(n40), .B0(n742), .B1(n605), .Y(n465) );
  OAI22XL U1183 ( .A0(n620), .A1(n33), .B0(n36), .B1(n621), .Y(n481) );
  OAI22XL U1184 ( .A0(n653), .A1(n24), .B0(n652), .B1(n21), .Y(n510) );
  NAND2X1 U1185 ( .A(n388), .B(n395), .Y(n169) );
  CMPR42X1 U1186 ( .A(n511), .B(n429), .C(n466), .D(n384), .ICI(n375), .S(n373), .ICO(n371), .CO(n372) );
  OAI22XL U1187 ( .A0(n607), .A1(n40), .B0(n42), .B1(n758), .Y(n429) );
  OAI22XL U1188 ( .A0(n606), .A1(n742), .B0(n605), .B1(n40), .Y(n466) );
  OAI22XL U1189 ( .A0(n654), .A1(n24), .B0(n653), .B1(n21), .Y(n511) );
  CMPR42X1 U1190 ( .A(n557), .B(n495), .C(n480), .D(n428), .ICI(n365), .S(n353), .ICO(n351), .CO(n352) );
  OAI22XL U1191 ( .A0(n589), .A1(n46), .B0(n48), .B1(n757), .Y(n428) );
  OAI22XL U1192 ( .A0(n620), .A1(n743), .B0(n619), .B1(n33), .Y(n480) );
  OAI22XL U1193 ( .A0(n636), .A1(n29), .B0(n635), .B1(n28), .Y(n495) );
  CMPR42X1 U1194 ( .A(n539), .B(n447), .C(n478), .D(n462), .ICI(n340), .S(n331), .ICO(n329), .CO(n330) );
  OAI22XL U1195 ( .A0(n602), .A1(n742), .B0(n601), .B1(n40), .Y(n462) );
  OAI22XL U1196 ( .A0(n618), .A1(n743), .B0(n617), .B1(n33), .Y(n478) );
  OAI22XL U1197 ( .A0(n586), .A1(n47), .B0(n45), .B1(n585), .Y(n447) );
  CMPR42X1 U1198 ( .A(n522), .B(n477), .C(n446), .D(n332), .ICI(n323), .S(n320), .ICO(n318), .CO(n319) );
  OAI22XL U1199 ( .A0(n584), .A1(n45), .B0(n47), .B1(n585), .Y(n446) );
  OAI22XL U1200 ( .A0(n617), .A1(n743), .B0(n616), .B1(n33), .Y(n477) );
  OAI22XL U1201 ( .A0(n664), .A1(n16), .B0(n665), .B1(n18), .Y(n522) );
  CMPR42X1 U1202 ( .A(n312), .B(n505), .C(n459), .D(n444), .ICI(n313), .S(n301), .ICO(n299), .CO(n300) );
  OAI22XL U1203 ( .A0(n583), .A1(n47), .B0(n582), .B1(n45), .Y(n444) );
  OAI22XL U1204 ( .A0(n599), .A1(n742), .B0(n598), .B1(n40), .Y(n459) );
  OAI22XL U1205 ( .A0(n646), .A1(n22), .B0(n647), .B1(n24), .Y(n505) );
  CLKINVX1 U1206 ( .A(n81), .Y(product_1_) );
  NAND2X1 U1207 ( .A(n427), .B(n553), .Y(n206) );
  CMPR42X1 U1208 ( .A(n562), .B(n485), .C(n546), .D(n514), .ICI(n530), .S(n399), .ICO(n397), .CO(n398) );
  OAI22XL U1209 ( .A0(n673), .A1(n746), .B0(n672), .B1(n15), .Y(n530) );
  OAI22XL U1210 ( .A0(n656), .A1(n21), .B0(n24), .B1(n657), .Y(n514) );
  NAND2X1 U1211 ( .A(n421), .B(n424), .Y(n198) );
  CMPR42X1 U1212 ( .A(n492), .B(n538), .C(n325), .D(n335), .ICI(n461), .S(n323), .ICO(n321), .CO(n322) );
  OAI22XL U1213 ( .A0(n601), .A1(n742), .B0(n600), .B1(n40), .Y(n461) );
  OAI22XL U1214 ( .A0(n12), .A1(n681), .B0(n680), .B1(n10), .Y(n538) );
  OR2X1 U1215 ( .A(n555), .B(n507), .Y(n335) );
  ADDHXL U1216 ( .A(n543), .B(n527), .CO(n376), .S(n377) );
  OAI22XL U1217 ( .A0(n12), .A1(n686), .B0(n685), .B1(n10), .Y(n543) );
  OAI22XL U1218 ( .A0(n670), .A1(n746), .B0(n669), .B1(n16), .Y(n527) );
  OAI22XL U1219 ( .A0(n674), .A1(n15), .B0(n746), .B1(n675), .Y(n532) );
  ADDFXL U1220 ( .A(n544), .B(n560), .CI(n392), .CO(n384), .S(n385) );
  OAI22XL U1221 ( .A0(n6), .A1(n703), .B0(n702), .B1(n3), .Y(n560) );
  OAI22XL U1222 ( .A0(n12), .A1(n687), .B0(n686), .B1(n10), .Y(n544) );
  ADDHXL U1223 ( .A(n551), .B(n567), .CO(n422), .S(n423) );
  OAI22XL U1224 ( .A0(n694), .A1(n747), .B0(n693), .B1(n9), .Y(n551) );
  OAI22XL U1225 ( .A0(n701), .A1(n3), .B0(n6), .B1(n702), .Y(n559) );
  OAI22XL U1226 ( .A0(n29), .A1(n631), .B0(n630), .B1(n28), .Y(n304) );
  OAI22XL U1227 ( .A0(n48), .A1(n579), .B0(n46), .B1(n578), .Y(n272) );
  CMPR42X1 U1228 ( .A(n504), .B(n299), .C(n293), .D(n300), .ICI(n296), .S(n290), .ICO(n288), .CO(n289) );
  OAI22XL U1229 ( .A0(n646), .A1(n24), .B0(n645), .B1(n22), .Y(n504) );
  CMPR42X1 U1230 ( .A(n489), .B(n291), .C(n285), .D(n292), .ICI(n288), .S(n282), .ICO(n280), .CO(n281) );
  OAI22XL U1231 ( .A0(n628), .A1(n28), .B0(n629), .B1(n744), .Y(n489) );
  CMPR42X1 U1232 ( .A(n454), .B(n270), .C(n266), .D(n470), .ICI(n267), .S(n264), .ICO(n262), .CO(n263) );
  OAI22XL U1233 ( .A0(n610), .A1(n36), .B0(n609), .B1(n34), .Y(n470) );
  OAI22XL U1234 ( .A0(n593), .A1(n40), .B0(n42), .B1(n594), .Y(n454) );
  CMPR42X1 U1235 ( .A(n472), .B(n283), .C(n279), .D(n284), .ICI(n280), .S(n276), .ICO(n274), .CO(n275) );
  OAI22XL U1236 ( .A0(n611), .A1(n34), .B0(n36), .B1(n612), .Y(n472) );
  CMPR42X1 U1237 ( .A(n277), .B(n271), .C(n471), .D(n278), .ICI(n274), .S(n269), .ICO(n267), .CO(n268) );
  OAI22XL U1238 ( .A0(n610), .A1(n34), .B0(n611), .B1(n36), .Y(n471) );
  OAI22XL U1239 ( .A0(n42), .A1(n596), .B0(n595), .B1(n40), .Y(n456) );
  OAI22XL U1240 ( .A0(n29), .A1(n632), .B0(n631), .B1(n28), .Y(n491) );
  CMPR42X1 U1241 ( .A(n458), .B(n490), .C(n302), .D(n295), .ICI(n443), .S(n293), .ICO(n291), .CO(n292) );
  OAI22XL U1242 ( .A0(n582), .A1(n47), .B0(n581), .B1(n45), .Y(n443) );
  OAI22XL U1243 ( .A0(n598), .A1(n742), .B0(n597), .B1(n40), .Y(n458) );
  OAI22XL U1244 ( .A0(n629), .A1(n28), .B0(n29), .B1(n630), .Y(n490) );
  CMPR42X1 U1245 ( .A(n286), .B(n456), .C(n503), .D(n441), .ICI(n488), .S(n279), .ICO(n277), .CO(n278) );
  OAI22XL U1246 ( .A0(n628), .A1(n744), .B0(n627), .B1(n28), .Y(n488) );
  OAI22XL U1247 ( .A0(n580), .A1(n47), .B0(n46), .B1(n579), .Y(n441) );
  CMPR42X1 U1248 ( .A(n457), .B(n473), .C(n287), .D(n294), .ICI(n442), .S(n285), .ICO(n283), .CO(n284) );
  OAI22XL U1249 ( .A0(n581), .A1(n47), .B0(n580), .B1(n45), .Y(n442) );
  OAI22XL U1250 ( .A0(n36), .A1(n613), .B0(n612), .B1(n34), .Y(n473) );
  OAI22XL U1251 ( .A0(n42), .A1(n597), .B0(n596), .B1(n40), .Y(n457) );
  ADDFXL U1252 ( .A(n455), .B(n487), .CI(n273), .CO(n270), .S(n271) );
  OAI22XL U1253 ( .A0(n42), .A1(n595), .B0(n594), .B1(n40), .Y(n455) );
  OAI22XL U1254 ( .A0(n744), .A1(n627), .B0(n626), .B1(n28), .Y(n487) );
  CLKINVX1 U1255 ( .A(n272), .Y(n273) );
  ADDFXL U1256 ( .A(n475), .B(n520), .CI(n305), .CO(n302), .S(n303) );
  OAI22XL U1257 ( .A0(n18), .A1(n663), .B0(n662), .B1(n16), .Y(n520) );
  OAI22XL U1258 ( .A0(n36), .A1(n615), .B0(n614), .B1(n34), .Y(n475) );
  CLKINVX1 U1259 ( .A(n304), .Y(n305) );
  ADDFXL U1260 ( .A(n272), .B(n440), .CI(n486), .CO(n265), .S(n266) );
  OAI22XL U1261 ( .A0(n48), .A1(n578), .B0(n46), .B1(n577), .Y(n440) );
  ADDFXL U1262 ( .A(n304), .B(n474), .CI(n519), .CO(n294), .S(n295) );
  OAI22XL U1263 ( .A0(n36), .A1(n614), .B0(n613), .B1(n34), .Y(n474) );
  CLKINVX1 U1264 ( .A(n43), .Y(n757) );
  OAI22XL U1265 ( .A0(n42), .A1(n591), .B0(n590), .B1(n40), .Y(n252) );
  OAI22XL U1266 ( .A0(n48), .A1(n577), .B0(n46), .B1(n576), .Y(n260) );
  CMPR42X1 U1267 ( .A(n260), .B(n468), .C(n439), .D(n452), .ICI(n257), .S(n256), .ICO(n254), .CO(n255) );
  OAI22XL U1268 ( .A0(n575), .A1(n46), .B0(n48), .B1(n576), .Y(n439) );
  OAI22XL U1269 ( .A0(n592), .A1(n42), .B0(n591), .B1(n40), .Y(n452) );
  CMPR42X1 U1270 ( .A(n469), .B(n261), .C(n265), .D(n453), .ICI(n262), .S(n259), .ICO(n257), .CO(n258) );
  OAI22XL U1271 ( .A0(n36), .A1(n609), .B0(n608), .B1(n34), .Y(n469) );
  OAI22XL U1272 ( .A0(n592), .A1(n40), .B0(n593), .B1(n42), .Y(n453) );
  CLKINVX1 U1273 ( .A(n260), .Y(n261) );
  OAI22XL U1274 ( .A0(n574), .A1(n48), .B0(n46), .B1(n573), .Y(n437) );
  CLKINVX1 U1275 ( .A(n252), .Y(n253) );
  OAI22XL U1276 ( .A0(n574), .A1(n46), .B0(n575), .B1(n48), .Y(n438) );
  XNOR2X1 U1277 ( .A(n717), .B(n43), .Y(n573) );
  XNOR2X1 U1278 ( .A(n716), .B(n43), .Y(n572) );
  OAI22X1 U1279 ( .A0(n696), .A1(n12), .B0(n695), .B1(n9), .Y(n553) );
  OAI22XL U1280 ( .A0(n643), .A1(n28), .B0(n744), .B1(n760), .Y(n431) );
  CLKINVX1 U1281 ( .A(n25), .Y(n760) );
  NAND2BX1 U1282 ( .AN(n49), .B(n25), .Y(n643) );
  CMPR42X1 U1283 ( .A(n513), .B(n430), .C(n394), .D(n398), .ICI(n391), .S(n388), .ICO(n386), .CO(n387) );
  OAI22XL U1284 ( .A0(n625), .A1(n34), .B0(n36), .B1(n759), .Y(n430) );
  OAI22XL U1285 ( .A0(n656), .A1(n24), .B0(n655), .B1(n21), .Y(n513) );
  CLKINVX1 U1286 ( .A(n31), .Y(n759) );
  XNOR2X1 U1287 ( .A(n7), .B(n722), .Y(n686) );
  XNOR2X1 U1288 ( .A(n1), .B(n722), .Y(n704) );
  XNOR2X1 U1289 ( .A(n1), .B(n717), .Y(n699) );
  XNOR2X1 U1290 ( .A(n1), .B(n721), .Y(n703) );
  XNOR2X1 U1291 ( .A(n7), .B(n721), .Y(n685) );
  XNOR2X1 U1292 ( .A(n19), .B(n721), .Y(n649) );
  XNOR2X1 U1293 ( .A(n7), .B(n723), .Y(n687) );
  XNOR2X1 U1294 ( .A(n1), .B(n723), .Y(n705) );
  XNOR2X1 U1295 ( .A(n13), .B(n723), .Y(n669) );
  XNOR2X1 U1296 ( .A(n1), .B(n720), .Y(n702) );
  XNOR2X1 U1297 ( .A(n19), .B(n720), .Y(n648) );
  XNOR2X1 U1298 ( .A(n1), .B(n731), .Y(n713) );
  XNOR2X1 U1299 ( .A(n25), .B(n731), .Y(n641) );
  XNOR2X1 U1300 ( .A(n13), .B(n729), .Y(n675) );
  XNOR2X1 U1301 ( .A(n728), .B(n7), .Y(n692) );
  XNOR2X1 U1302 ( .A(n730), .B(n13), .Y(n676) );
  XNOR2X1 U1303 ( .A(n718), .B(n1), .Y(n700) );
  XNOR2X1 U1304 ( .A(n725), .B(n7), .Y(n689) );
  XNOR2X1 U1305 ( .A(n726), .B(n7), .Y(n690) );
  XNOR2X1 U1306 ( .A(n724), .B(n1), .Y(n706) );
  XNOR2X1 U1307 ( .A(n719), .B(n1), .Y(n701) );
  XNOR2X1 U1308 ( .A(n727), .B(n7), .Y(n691) );
  XNOR2X1 U1309 ( .A(n726), .B(n1), .Y(n708) );
  XNOR2X1 U1310 ( .A(n1), .B(n716), .Y(n698) );
  ADDHX1 U1311 ( .A(n569), .B(n434), .CO(n426), .S(n427) );
  ADDFX2 U1312 ( .A(n433), .B(n535), .CI(n423), .CO(n420), .S(n421) );
  OAI22XL U1313 ( .A0(n679), .A1(n16), .B0(n18), .B1(n762), .Y(n433) );
  OAI22XL U1314 ( .A0(n678), .A1(n746), .B0(n677), .B1(n15), .Y(n535) );
  CLKINVX1 U1315 ( .A(n13), .Y(n762) );
  CLKBUFX3 U1316 ( .A(n749), .Y(n46) );
  CLKBUFX3 U1317 ( .A(n754), .Y(n16) );
  CLKBUFX3 U1318 ( .A(n753), .Y(n22) );
  CLKBUFX3 U1319 ( .A(n752), .Y(n28) );
  CLKBUFX3 U1320 ( .A(n750), .Y(n40) );
  CLKBUFX3 U1321 ( .A(n751), .Y(n34) );
  CLKBUFX3 U1322 ( .A(n755), .Y(n10) );
  CLKBUFX3 U1323 ( .A(n749), .Y(n45) );
  CLKBUFX3 U1324 ( .A(n754), .Y(n15) );
  CLKBUFX3 U1325 ( .A(n753), .Y(n21) );
  CLKBUFX3 U1326 ( .A(n751), .Y(n33) );
  CLKBUFX3 U1327 ( .A(n755), .Y(n9) );
  CLKBUFX3 U1328 ( .A(n741), .Y(n47) );
  CLKBUFX3 U1329 ( .A(n756), .Y(n3) );
  CLKBUFX3 U1330 ( .A(n741), .Y(n48) );
  CLKBUFX3 U1331 ( .A(n746), .Y(n18) );
  CLKINVX1 U1332 ( .A(n19), .Y(n761) );
  CLKINVX1 U1333 ( .A(n37), .Y(n758) );
  XNOR2X1 U1334 ( .A(n19), .B(n717), .Y(n645) );
  XNOR2X1 U1335 ( .A(n19), .B(n716), .Y(n644) );
  XOR2X1 U1336 ( .A(a_5_), .B(a_4_), .Y(n738) );
  NAND2X1 U1337 ( .A(n737), .B(n753), .Y(n745) );
  XOR2X1 U1338 ( .A(a_7_), .B(a_6_), .Y(n737) );
  NAND2X1 U1339 ( .A(n736), .B(n752), .Y(n744) );
  XOR2X1 U1340 ( .A(a_9_), .B(a_8_), .Y(n736) );
  NAND2X1 U1341 ( .A(n735), .B(n751), .Y(n743) );
  XOR2X1 U1342 ( .A(a_11_), .B(a_10_), .Y(n735) );
  XOR2X1 U1343 ( .A(a_13_), .B(a_12_), .Y(n734) );
  XOR2X1 U1344 ( .A(a_3_), .B(a_2_), .Y(n739) );
  XOR2X1 U1345 ( .A(a_14_), .B(a_15_), .Y(n733) );
  NAND2X1 U1346 ( .A(n740), .B(n756), .Y(n748) );
  XOR2X1 U1347 ( .A(a_0_), .B(a_1_), .Y(n740) );
endmodule


module FFT_ultrafast2_shift_DW_mult_uns_10 ( a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_, 
        b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, product_31_, product_30_, 
        product_29_, product_28_, product_27_, product_26_, product_25_, 
        product_24_, product_23_, product_22_, product_21_, product_20_, 
        product_19_, product_18_, product_17_, product_16_, product_15_, 
        product_14_, product_13_, product_12_, product_11_, product_10_, 
        product_9_, product_8_, product_7_, product_6_, product_5_, product_4_, 
        product_3_, product_2_, product_1_, product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_, b_16_, b_15_, b_14_, b_13_, b_12_,
         b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_,
         b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n4, n5, n7, n13, n16, n17, n19, n21, n22, n24, n25, n28, n29, n31,
         n33, n34, n36, n37, n40, n41, n42, n43, n46, n48, n49, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n83, n86, n88, n89, n90, n91, n92, n94, n96, n97, n98, n99, n100,
         n102, n104, n105, n106, n107, n108, n110, n112, n113, n114, n115,
         n116, n118, n120, n121, n122, n123, n124, n126, n128, n129, n130,
         n131, n132, n134, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n164, n165, n166,
         n167, n168, n169, n171, n173, n174, n176, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n193,
         n195, n196, n198, n200, n201, n202, n204, n206, n207, n208, n209,
         n210, n212, n214, n215, n216, n217, n218, n219, n222, n224, n226,
         n228, n230, n232, n234, n235, n236, n238, n239, n242, n243, n247,
         n249, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n728, n729, n731, n733, n734, n735,
         n736, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857;

  OAI22X1 U699 ( .A0(n660), .A1(n24), .B0(n659), .B1(n21), .Y(n517) );
  OAI21X2 U700 ( .A0(n190), .A1(n202), .B0(n191), .Y(n189) );
  AOI21X4 U701 ( .A0(n157), .A1(n148), .B0(n149), .Y(n147) );
  OAI21X1 U702 ( .A0(n150), .A1(n156), .B0(n151), .Y(n149) );
  OAI22X1 U703 ( .A0(n643), .A1(n29), .B0(n642), .B1(n28), .Y(n500) );
  BUFX4 U704 ( .A(b_2_), .Y(n735) );
  AOI21X2 U705 ( .A0(n179), .A1(n841), .B0(n176), .Y(n174) );
  INVX1 U706 ( .A(n180), .Y(n179) );
  OAI21X2 U707 ( .A0(n180), .A1(n168), .B0(n169), .Y(n167) );
  AOI21X2 U708 ( .A0(n181), .A1(n189), .B0(n182), .Y(n180) );
  ADDHX1 U709 ( .A(n439), .B(n558), .CO(n431), .S(n432) );
  XNOR2X4 U710 ( .A(n185), .B(n73), .Y(product_9_) );
  OAI21X1 U711 ( .A0(n188), .A1(n186), .B0(n187), .Y(n185) );
  XNOR2X4 U712 ( .A(n735), .B(n1), .Y(n717) );
  ADDFHX2 U713 ( .A(n541), .B(n557), .CI(n573), .CO(n429), .S(n430) );
  OAI22X1 U714 ( .A0(n695), .A1(n760), .B0(n752), .B1(n700), .Y(n557) );
  OAI22X2 U715 ( .A0(n695), .A1(n752), .B0(n695), .B1(n760), .Y(n553) );
  ADDFHX2 U716 ( .A(n536), .B(n504), .CI(n411), .CO(n408), .S(n409) );
  OAI22X1 U717 ( .A0(n679), .A1(n17), .B0(n678), .B1(n759), .Y(n536) );
  OAI22X1 U718 ( .A0(n659), .A1(n750), .B0(n658), .B1(n21), .Y(n516) );
  OAI22X1 U719 ( .A0(n665), .A1(n750), .B0(n664), .B1(n21), .Y(n522) );
  BUFX12 U720 ( .A(n750), .Y(n24) );
  OAI22X4 U721 ( .A0(n663), .A1(n21), .B0(n750), .B1(n664), .Y(n521) );
  NAND2X4 U722 ( .A(n742), .B(n758), .Y(n750) );
  OAI21X4 U723 ( .A0(n138), .A1(n158), .B0(n139), .Y(n137) );
  AOI21X2 U724 ( .A0(n167), .A1(n159), .B0(n160), .Y(n158) );
  AOI21X1 U725 ( .A0(n140), .A1(n149), .B0(n141), .Y(n139) );
  OAI21X4 U726 ( .A0(n116), .A1(n114), .B0(n115), .Y(n113) );
  AOI21X4 U727 ( .A0(n121), .A1(n846), .B0(n118), .Y(n116) );
  INVXL U728 ( .A(n19), .Y(n766) );
  OAI22X1 U729 ( .A0(n684), .A1(n16), .B0(n17), .B1(n767), .Y(n438) );
  XNOR2X2 U730 ( .A(n19), .B(n736), .Y(n664) );
  XNOR2X1 U731 ( .A(n731), .B(n19), .Y(n659) );
  OAI22XL U732 ( .A0(n720), .A1(n4), .B0(n753), .B1(n852), .Y(n440) );
  NAND2BX1 U733 ( .AN(n49), .B(n1), .Y(n720) );
  OAI22XL U734 ( .A0(n716), .A1(n4), .B0(n717), .B1(n5), .Y(n574) );
  OAI22XL U735 ( .A0(n701), .A1(n752), .B0(n700), .B1(n760), .Y(n558) );
  OAI22XL U736 ( .A0(n702), .A1(n760), .B0(n752), .B1(n768), .Y(n439) );
  XNOR2X1 U737 ( .A(n7), .B(n736), .Y(n700) );
  NAND2X1 U738 ( .A(n432), .B(n574), .Y(n214) );
  OR2X1 U739 ( .A(n432), .B(n574), .Y(n844) );
  XNOR2X1 U740 ( .A(n49), .B(n19), .Y(n665) );
  XNOR2X1 U741 ( .A(n735), .B(n13), .Y(n681) );
  XNOR2X1 U742 ( .A(n734), .B(n13), .Y(n680) );
  OAI22XL U743 ( .A0(n666), .A1(n22), .B0(n24), .B1(n766), .Y(n437) );
  NAND2BX1 U744 ( .AN(n49), .B(n19), .Y(n666) );
  OAI22XL U745 ( .A0(n717), .A1(n5), .B0(n714), .B1(n4), .Y(n572) );
  CMPR42X1 U746 ( .A(n435), .B(n486), .C(n398), .D(n502), .ICI(n402), .S(n396), 
        .ICO(n394), .CO(n395) );
  XNOR2X1 U747 ( .A(n13), .B(n729), .Y(n675) );
  XNOR2X1 U748 ( .A(n7), .B(n724), .Y(n688) );
  OAI21XL U749 ( .A0(n183), .A1(n187), .B0(n184), .Y(n182) );
  OR2X1 U750 ( .A(n419), .B(n423), .Y(n842) );
  CLKINVX1 U751 ( .A(n178), .Y(n176) );
  CMPR42X1 U752 ( .A(n500), .B(n470), .C(n389), .D(n484), .ICI(n386), .S(n378), 
        .ICO(n376), .CO(n377) );
  OAI22XL U753 ( .A0(n611), .A1(n41), .B0(n610), .B1(n40), .Y(n470) );
  ADDFXL U754 ( .A(n382), .B(n516), .CI(n434), .CO(n379), .S(n380) );
  CLKBUFX3 U755 ( .A(a_1_), .Y(n1) );
  CLKBUFX3 U756 ( .A(a_7_), .Y(n19) );
  XNOR2X1 U757 ( .A(a_5_), .B(a_6_), .Y(n758) );
  CLKBUFX3 U758 ( .A(a_5_), .Y(n13) );
  CLKINVX1 U759 ( .A(n183), .Y(n242) );
  OA21XL U760 ( .A0(n166), .A1(n164), .B0(n165), .Y(n855) );
  OAI22X1 U761 ( .A0(n577), .A1(n46), .B0(n48), .B1(n578), .Y(n251) );
  AOI21X1 U762 ( .A0(n113), .A1(n847), .B0(n110), .Y(n108) );
  OAI21X1 U763 ( .A0(n108), .A1(n106), .B0(n107), .Y(n105) );
  AOI21X1 U764 ( .A0(n97), .A1(n848), .B0(n94), .Y(n92) );
  AOI21X1 U765 ( .A0(n129), .A1(n843), .B0(n126), .Y(n124) );
  CLKINVX1 U766 ( .A(n128), .Y(n126) );
  OAI21X1 U767 ( .A0(n132), .A1(n130), .B0(n131), .Y(n129) );
  CLKINVX1 U768 ( .A(n120), .Y(n118) );
  CLKBUFX3 U769 ( .A(b_3_), .Y(n734) );
  CLKBUFX3 U770 ( .A(b_9_), .Y(n728) );
  OR2X1 U771 ( .A(n393), .B(n400), .Y(n838) );
  OR2X1 U772 ( .A(n424), .B(n425), .Y(n839) );
  CLKBUFX3 U773 ( .A(n746), .Y(n48) );
  OR2X1 U774 ( .A(n322), .B(n332), .Y(n840) );
  OR2X1 U775 ( .A(n401), .B(n406), .Y(n841) );
  OR2X1 U776 ( .A(n312), .B(n303), .Y(n843) );
  OR2X1 U777 ( .A(n426), .B(n429), .Y(n845) );
  OR2X1 U778 ( .A(n294), .B(n287), .Y(n846) );
  OR2X1 U779 ( .A(n274), .B(n280), .Y(n847) );
  OR2X1 U780 ( .A(n256), .B(n260), .Y(n848) );
  OR2X1 U781 ( .A(n268), .B(n264), .Y(n849) );
  OR2X1 U782 ( .A(n253), .B(n252), .Y(n850) );
  NAND2X1 U783 ( .A(n741), .B(n757), .Y(n749) );
  BUFX4 U784 ( .A(n749), .Y(n29) );
  BUFX4 U785 ( .A(n751), .Y(n17) );
  XNOR2X1 U786 ( .A(a_7_), .B(a_8_), .Y(n757) );
  BUFX4 U787 ( .A(n757), .Y(n28) );
  OAI21X1 U788 ( .A0(n147), .A1(n145), .B0(n146), .Y(n144) );
  XNOR2X2 U789 ( .A(a_3_), .B(a_4_), .Y(n759) );
  CLKBUFX3 U790 ( .A(n758), .Y(n21) );
  ADDHX2 U791 ( .A(n438), .B(n540), .CO(n427), .S(n428) );
  CLKBUFX6 U792 ( .A(a_3_), .Y(n7) );
  XNOR2X4 U793 ( .A(n731), .B(n7), .Y(n695) );
  XNOR2X1 U794 ( .A(n735), .B(n31), .Y(n627) );
  OAI22X1 U795 ( .A0(n716), .A1(n5), .B0(n717), .B1(n4), .Y(n573) );
  CMPR42X2 U796 ( .A(n523), .B(n539), .C(n571), .D(n555), .ICI(n427), .S(n424), 
        .ICO(n422), .CO(n423) );
  OAI22X1 U797 ( .A0(n681), .A1(n759), .B0(n17), .B1(n682), .Y(n539) );
  NOR2X2 U798 ( .A(n407), .B(n413), .Y(n183) );
  OAI22X1 U799 ( .A0(n752), .A1(n694), .B0(n693), .B1(n760), .Y(n551) );
  XNOR2X1 U800 ( .A(n7), .B(n729), .Y(n693) );
  XNOR2X4 U801 ( .A(n728), .B(n7), .Y(n692) );
  CMPR32X2 U802 ( .A(n572), .B(n556), .C(n428), .CO(n425), .S(n426) );
  ADDHX1 U803 ( .A(n570), .B(n437), .CO(n420), .S(n421) );
  ADDHX1 U804 ( .A(n566), .B(n534), .CO(n397), .S(n398) );
  OAI22X1 U805 ( .A0(n17), .A1(n676), .B0(n675), .B1(n16), .Y(n533) );
  OAI22X1 U806 ( .A0(n678), .A1(n17), .B0(n676), .B1(n16), .Y(n534) );
  BUFX20 U807 ( .A(a_9_), .Y(n25) );
  XNOR2X1 U808 ( .A(n49), .B(n7), .Y(n701) );
  NAND2BX1 U809 ( .AN(n49), .B(n7), .Y(n702) );
  NAND2BX1 U810 ( .AN(n49), .B(n13), .Y(n684) );
  XNOR2XL U811 ( .A(n49), .B(n25), .Y(n647) );
  BUFX20 U812 ( .A(b_0_), .Y(n49) );
  OAI22X1 U813 ( .A0(n683), .A1(n17), .B0(n682), .B1(n759), .Y(n540) );
  XNOR2X4 U814 ( .A(a_1_), .B(a_2_), .Y(n760) );
  XOR2XL U815 ( .A(a_5_), .B(a_4_), .Y(n743) );
  NAND2X1 U816 ( .A(n731), .B(n1), .Y(n853) );
  NAND2X2 U817 ( .A(n851), .B(n852), .Y(n854) );
  NAND2X4 U818 ( .A(n853), .B(n854), .Y(n713) );
  INVX1 U819 ( .A(n731), .Y(n851) );
  INVXL U820 ( .A(n1), .Y(n852) );
  OAI22X1 U821 ( .A0(n713), .A1(n5), .B0(n712), .B1(n4), .Y(n570) );
  OAI22X1 U822 ( .A0(n714), .A1(n5), .B0(n713), .B1(n4), .Y(n571) );
  XOR2X1 U823 ( .A(n116), .B(n59), .Y(product_23_) );
  INVX1 U824 ( .A(n173), .Y(n171) );
  INVX1 U825 ( .A(n200), .Y(n198) );
  XOR2XL U826 ( .A(n124), .B(n61), .Y(product_21_) );
  NAND2X1 U827 ( .A(n840), .B(n136), .Y(n64) );
  BUFX4 U828 ( .A(n753), .Y(n5) );
  CLKBUFX3 U829 ( .A(a_15_), .Y(n43) );
  OAI22XL U830 ( .A0(n17), .A1(n671), .B0(n670), .B1(n16), .Y(n528) );
  XNOR2XL U831 ( .A(n7), .B(b_12_), .Y(n689) );
  CLKBUFX3 U832 ( .A(a_11_), .Y(n31) );
  XNOR2X1 U833 ( .A(n723), .B(n7), .Y(n687) );
  INVX1 U834 ( .A(n202), .Y(n201) );
  NAND2XL U835 ( .A(n140), .B(n148), .Y(n138) );
  XNOR2XL U836 ( .A(b_7_), .B(n13), .Y(n676) );
  OAI22X1 U837 ( .A0(n630), .A1(n34), .B0(n36), .B1(n764), .Y(n435) );
  OAI22X1 U838 ( .A0(n629), .A1(n36), .B0(n628), .B1(n33), .Y(n486) );
  XNOR2XL U839 ( .A(n733), .B(n31), .Y(n625) );
  XNOR2XL U840 ( .A(n728), .B(n19), .Y(n656) );
  XNOR2XL U841 ( .A(n734), .B(n37), .Y(n608) );
  XNOR2XL U842 ( .A(n25), .B(n729), .Y(n639) );
  XNOR2XL U843 ( .A(b_7_), .B(n25), .Y(n640) );
  XNOR2XL U844 ( .A(n728), .B(n13), .Y(n674) );
  CLKBUFX3 U845 ( .A(a_13_), .Y(n37) );
  XOR2X1 U846 ( .A(n166), .B(n70), .Y(product_12_) );
  INVXL U847 ( .A(n164), .Y(n239) );
  INVXL U848 ( .A(n142), .Y(n234) );
  INVXL U849 ( .A(n150), .Y(n236) );
  OAI21XL U850 ( .A0(n142), .A1(n146), .B0(n143), .Y(n141) );
  INVXL U851 ( .A(n114), .Y(n228) );
  INVXL U852 ( .A(n122), .Y(n230) );
  OAI21X1 U853 ( .A0(n208), .A1(n210), .B0(n209), .Y(n207) );
  NAND2X1 U854 ( .A(n385), .B(n392), .Y(n165) );
  INVXL U855 ( .A(n216), .Y(n249) );
  NAND2X1 U856 ( .A(n576), .B(n440), .Y(n219) );
  CMPR42X1 U857 ( .A(n518), .B(n550), .C(n403), .D(n399), .ICI(n396), .S(n393), 
        .ICO(n391), .CO(n392) );
  AO21XL U858 ( .A0(n42), .A1(n40), .B0(n595), .Y(n456) );
  XNOR2X1 U859 ( .A(b_7_), .B(n1), .Y(n712) );
  XNOR2X1 U860 ( .A(n7), .B(n722), .Y(n686) );
  OAI22X1 U861 ( .A0(n648), .A1(n28), .B0(n29), .B1(n765), .Y(n436) );
  CLKBUFX2 U862 ( .A(n747), .Y(n42) );
  NAND2X2 U863 ( .A(n740), .B(n756), .Y(n748) );
  INVX3 U864 ( .A(n158), .Y(n157) );
  XOR2X1 U865 ( .A(n855), .B(n69), .Y(product_13_) );
  NAND2XL U866 ( .A(n236), .B(n151), .Y(n67) );
  XNOR2XL U867 ( .A(n157), .B(n68), .Y(product_14_) );
  NAND2XL U868 ( .A(n153), .B(n156), .Y(n68) );
  INVXL U869 ( .A(n156), .Y(n154) );
  XOR2XL U870 ( .A(n108), .B(n57), .Y(product_25_) );
  XOR2XL U871 ( .A(n78), .B(n210), .Y(product_4_) );
  NAND2XL U872 ( .A(n247), .B(n209), .Y(n78) );
  XNOR2XL U873 ( .A(n79), .B(n215), .Y(product_3_) );
  NAND2XL U874 ( .A(n844), .B(n214), .Y(n79) );
  NAND2XL U875 ( .A(n249), .B(n217), .Y(n80) );
  XOR2XL U876 ( .A(n188), .B(n74), .Y(product_8_) );
  NAND2XL U877 ( .A(n243), .B(n187), .Y(n74) );
  NAND2XL U878 ( .A(n842), .B(n195), .Y(n75) );
  OAI21X4 U879 ( .A0(n100), .A1(n98), .B0(n99), .Y(n97) );
  XNOR2XL U880 ( .A(n207), .B(n77), .Y(product_5_) );
  NAND2XL U881 ( .A(n845), .B(n206), .Y(n77) );
  XNOR2X1 U882 ( .A(n856), .B(n51), .Y(product_31_) );
  AO21XL U883 ( .A0(n89), .A1(n850), .B0(n86), .Y(n856) );
  NOR2X1 U884 ( .A(n355), .B(n365), .Y(n150) );
  NOR2X1 U885 ( .A(n366), .B(n374), .Y(n155) );
  NOR2X1 U886 ( .A(n385), .B(n392), .Y(n164) );
  XOR2XL U887 ( .A(n100), .B(n55), .Y(product_27_) );
  CLKBUFX2 U888 ( .A(b_14_), .Y(n723) );
  NOR2X1 U889 ( .A(n333), .B(n343), .Y(n142) );
  NOR2X1 U890 ( .A(n344), .B(n354), .Y(n145) );
  NOR2X1 U891 ( .A(n313), .B(n321), .Y(n130) );
  NOR2X1 U892 ( .A(n302), .B(n295), .Y(n122) );
  NOR2X1 U893 ( .A(n281), .B(n286), .Y(n114) );
  NOR2X1 U894 ( .A(n269), .B(n273), .Y(n106) );
  NOR2X1 U895 ( .A(n254), .B(n255), .Y(n90) );
  CMPR42X2 U896 ( .A(n415), .B(n520), .C(n568), .D(n409), .ICI(n412), .S(n407), 
        .ICO(n405), .CO(n406) );
  NOR2BXL U897 ( .AN(n49), .B(n760), .Y(n559) );
  CLKBUFX2 U898 ( .A(b_8_), .Y(n729) );
  NOR2BXL U899 ( .AN(n49), .B(n33), .Y(n487) );
  NOR2X1 U900 ( .A(n414), .B(n418), .Y(n186) );
  NOR2X1 U901 ( .A(n575), .B(n559), .Y(n216) );
  NOR2X1 U902 ( .A(n430), .B(n431), .Y(n208) );
  NAND2BXL U903 ( .AN(n218), .B(n219), .Y(n81) );
  NOR2XL U904 ( .A(n576), .B(n440), .Y(n218) );
  XNOR2XL U905 ( .A(n735), .B(n43), .Y(n591) );
  XNOR2XL U906 ( .A(n734), .B(n43), .Y(n590) );
  XNOR2XL U907 ( .A(n49), .B(n43), .Y(n593) );
  NOR2BXL U908 ( .AN(n49), .B(n4), .Y(product_0_) );
  NAND2BXL U909 ( .AN(n49), .B(n43), .Y(n594) );
  XNOR2XL U910 ( .A(n733), .B(n43), .Y(n589) );
  XNOR2XL U911 ( .A(n733), .B(n43), .Y(n588) );
  XNOR2XL U912 ( .A(n731), .B(n43), .Y(n587) );
  XNOR2XL U913 ( .A(b_7_), .B(n43), .Y(n586) );
  XNOR2XL U914 ( .A(n728), .B(n43), .Y(n584) );
  XNOR2XL U915 ( .A(n729), .B(n43), .Y(n585) );
  OAI22XL U916 ( .A0(n748), .A1(n622), .B0(n621), .B1(n33), .Y(n329) );
  AO21XL U917 ( .A0(n749), .A1(n28), .B0(n631), .Y(n488) );
  XNOR2XL U918 ( .A(b_11_), .B(n43), .Y(n582) );
  XNOR2XL U919 ( .A(b_12_), .B(n43), .Y(n581) );
  XNOR2XL U920 ( .A(n43), .B(n722), .Y(n583) );
  NOR2X1 U921 ( .A(n261), .B(n263), .Y(n98) );
  ADDFXL U922 ( .A(n258), .B(n259), .CI(n457), .CO(n255), .S(n256) );
  XNOR2XL U923 ( .A(n723), .B(n43), .Y(n579) );
  ADDFXL U924 ( .A(n442), .B(n257), .CI(n456), .CO(n253), .S(n254) );
  AO21XL U925 ( .A0(n48), .A1(n46), .B0(n577), .Y(n441) );
  ADDHX1 U926 ( .A(n552), .B(n436), .CO(n410), .S(n411) );
  OAI22X1 U927 ( .A0(n695), .A1(n752), .B0(n694), .B1(n760), .Y(n552) );
  XNOR2XL U928 ( .A(b_5_), .B(n1), .Y(n714) );
  XNOR2XL U929 ( .A(n735), .B(n25), .Y(n645) );
  XNOR2XL U930 ( .A(b_5_), .B(n19), .Y(n660) );
  XNOR2XL U931 ( .A(b_5_), .B(n25), .Y(n642) );
  XNOR2XL U932 ( .A(n733), .B(n19), .Y(n661) );
  XNOR2XL U933 ( .A(n733), .B(n25), .Y(n643) );
  XNOR2XL U934 ( .A(n734), .B(n19), .Y(n662) );
  XNOR2XL U935 ( .A(n734), .B(n25), .Y(n644) );
  XNOR2XL U936 ( .A(n734), .B(n31), .Y(n626) );
  CLKBUFX2 U937 ( .A(n758), .Y(n22) );
  XNOR2XL U938 ( .A(n49), .B(n13), .Y(n683) );
  XNOR2XL U939 ( .A(n49), .B(n31), .Y(n629) );
  XNOR2XL U940 ( .A(n49), .B(n37), .Y(n611) );
  NAND2BXL U941 ( .AN(n49), .B(n25), .Y(n648) );
  NAND2BXL U942 ( .AN(n49), .B(n31), .Y(n630) );
  NAND2BXL U943 ( .AN(n49), .B(n37), .Y(n612) );
  NOR2BXL U944 ( .AN(n49), .B(n16), .Y(n541) );
  XNOR2XL U945 ( .A(n13), .B(b_12_), .Y(n671) );
  XNOR2XL U946 ( .A(b_7_), .B(n19), .Y(n658) );
  XNOR2XL U947 ( .A(n735), .B(n37), .Y(n609) );
  XNOR2XL U948 ( .A(n731), .B(n25), .Y(n641) );
  XNOR2XL U949 ( .A(n731), .B(n31), .Y(n623) );
  XNOR2XL U950 ( .A(n733), .B(n37), .Y(n607) );
  XNOR2XL U951 ( .A(n733), .B(n37), .Y(n606) );
  XNOR2XL U952 ( .A(n728), .B(n25), .Y(n638) );
  XNOR2XL U953 ( .A(b_11_), .B(n13), .Y(n672) );
  XNOR2XL U954 ( .A(b_11_), .B(n19), .Y(n654) );
  XNOR2XL U955 ( .A(n19), .B(b_12_), .Y(n653) );
  XNOR2XL U956 ( .A(n721), .B(n7), .Y(n685) );
  XNOR2XL U957 ( .A(n19), .B(n729), .Y(n657) );
  XNOR2XL U958 ( .A(n13), .B(n722), .Y(n673) );
  XNOR2XL U959 ( .A(n19), .B(n722), .Y(n655) );
  CLKBUFX2 U960 ( .A(n755), .Y(n40) );
  XNOR2XL U961 ( .A(n723), .B(n31), .Y(n615) );
  XNOR2XL U962 ( .A(n31), .B(n729), .Y(n621) );
  XNOR2XL U963 ( .A(n723), .B(n13), .Y(n669) );
  XNOR2XL U964 ( .A(b_7_), .B(n37), .Y(n604) );
  XNOR2XL U965 ( .A(n723), .B(n19), .Y(n651) );
  XNOR2XL U966 ( .A(n723), .B(n25), .Y(n633) );
  XNOR2XL U967 ( .A(n731), .B(n37), .Y(n605) );
  XNOR2XL U968 ( .A(n728), .B(n31), .Y(n620) );
  XNOR2XL U969 ( .A(b_11_), .B(n25), .Y(n636) );
  XNOR2XL U970 ( .A(n728), .B(n37), .Y(n602) );
  XNOR2XL U971 ( .A(b_11_), .B(n31), .Y(n618) );
  XNOR2XL U972 ( .A(b_11_), .B(n37), .Y(n600) );
  XNOR2XL U973 ( .A(n25), .B(b_12_), .Y(n635) );
  XNOR2XL U974 ( .A(n31), .B(b_12_), .Y(n617) );
  XNOR2XL U975 ( .A(n37), .B(b_12_), .Y(n599) );
  XNOR2XL U976 ( .A(n721), .B(n13), .Y(n667) );
  XNOR2XL U977 ( .A(n721), .B(n19), .Y(n649) );
  XNOR2XL U978 ( .A(n721), .B(n25), .Y(n631) );
  XNOR2XL U979 ( .A(n37), .B(n729), .Y(n603) );
  XNOR2XL U980 ( .A(n13), .B(n722), .Y(n668) );
  XNOR2XL U981 ( .A(n25), .B(n722), .Y(n637) );
  XNOR2XL U982 ( .A(n31), .B(n722), .Y(n619) );
  XNOR2XL U983 ( .A(n19), .B(n722), .Y(n650) );
  XNOR2XL U984 ( .A(n25), .B(n722), .Y(n632) );
  OAI22XL U985 ( .A0(n36), .A1(n616), .B0(n615), .B1(n34), .Y(n277) );
  XNOR2XL U986 ( .A(n721), .B(n31), .Y(n613) );
  XNOR2XL U987 ( .A(n721), .B(n37), .Y(n595) );
  XNOR2XL U988 ( .A(n37), .B(n722), .Y(n601) );
  XNOR2XL U989 ( .A(n31), .B(n722), .Y(n614) );
  OAI22XL U990 ( .A0(n42), .A1(n598), .B0(n597), .B1(n40), .Y(n265) );
  AO21XL U991 ( .A0(n36), .A1(n34), .B0(n613), .Y(n472) );
  XNOR2XL U992 ( .A(n723), .B(n37), .Y(n597) );
  XNOR2XL U993 ( .A(n37), .B(n722), .Y(n596) );
  OAI22XL U994 ( .A0(n579), .A1(n46), .B0(n48), .B1(n580), .Y(n257) );
  XNOR2X1 U995 ( .A(a_9_), .B(a_10_), .Y(n756) );
  NAND2X4 U996 ( .A(n744), .B(n760), .Y(n752) );
  INVX1 U997 ( .A(a_0_), .Y(n761) );
  XNOR2XL U998 ( .A(n13), .B(n724), .Y(n670) );
  XNOR2X1 U999 ( .A(a_13_), .B(a_14_), .Y(n754) );
  XNOR2XL U1000 ( .A(n19), .B(n724), .Y(n652) );
  XNOR2XL U1001 ( .A(n25), .B(n724), .Y(n634) );
  XNOR2XL U1002 ( .A(n43), .B(n724), .Y(n580) );
  CLKBUFX2 U1003 ( .A(b_1_), .Y(n736) );
  CLKBUFX2 U1004 ( .A(b_13_), .Y(n724) );
  CLKINVX1 U1005 ( .A(n167), .Y(n166) );
  XNOR2X1 U1006 ( .A(n179), .B(n72), .Y(product_10_) );
  NAND2X1 U1007 ( .A(n841), .B(n178), .Y(n72) );
  XNOR2X1 U1008 ( .A(n144), .B(n65), .Y(product_17_) );
  NAND2X1 U1009 ( .A(n234), .B(n143), .Y(n65) );
  NAND2X1 U1010 ( .A(n238), .B(n162), .Y(n69) );
  CLKINVX1 U1011 ( .A(n161), .Y(n238) );
  XNOR2X1 U1012 ( .A(n89), .B(n52), .Y(product_30_) );
  NAND2X1 U1013 ( .A(n850), .B(n88), .Y(n52) );
  XNOR2X1 U1014 ( .A(n105), .B(n56), .Y(product_26_) );
  NAND2X1 U1015 ( .A(n849), .B(n104), .Y(n56) );
  XNOR2X1 U1016 ( .A(n113), .B(n58), .Y(product_24_) );
  NAND2X1 U1017 ( .A(n847), .B(n112), .Y(n58) );
  XNOR2X1 U1018 ( .A(n121), .B(n60), .Y(product_22_) );
  NAND2X1 U1019 ( .A(n846), .B(n120), .Y(n60) );
  XNOR2X1 U1020 ( .A(n129), .B(n62), .Y(product_20_) );
  NAND2X1 U1021 ( .A(n843), .B(n128), .Y(n62) );
  XNOR2X1 U1022 ( .A(n137), .B(n64), .Y(product_18_) );
  NAND2X1 U1023 ( .A(n838), .B(n841), .Y(n168) );
  AOI21X1 U1024 ( .A0(n838), .A1(n176), .B0(n171), .Y(n169) );
  OAI21XL U1025 ( .A0(n161), .A1(n165), .B0(n162), .Y(n160) );
  NOR2X1 U1026 ( .A(n164), .B(n161), .Y(n159) );
  AOI21X1 U1027 ( .A0(n137), .A1(n840), .B0(n134), .Y(n132) );
  CLKINVX1 U1028 ( .A(n136), .Y(n134) );
  CLKINVX1 U1029 ( .A(n112), .Y(n110) );
  AOI21X1 U1030 ( .A0(n105), .A1(n849), .B0(n102), .Y(n100) );
  CLKINVX1 U1031 ( .A(n104), .Y(n102) );
  OAI21X1 U1032 ( .A0(n124), .A1(n122), .B0(n123), .Y(n121) );
  OAI21XL U1033 ( .A0(n92), .A1(n90), .B0(n91), .Y(n89) );
  NOR2X1 U1034 ( .A(n142), .B(n145), .Y(n140) );
  CLKBUFX3 U1035 ( .A(b_4_), .Y(n733) );
  CLKBUFX3 U1036 ( .A(b_6_), .Y(n731) );
  NOR2X1 U1037 ( .A(n155), .B(n150), .Y(n148) );
  XOR2X1 U1038 ( .A(n174), .B(n71), .Y(product_11_) );
  NAND2X1 U1039 ( .A(n838), .B(n173), .Y(n71) );
  XOR2X1 U1040 ( .A(n152), .B(n67), .Y(product_15_) );
  AOI21X1 U1041 ( .A0(n157), .A1(n153), .B0(n154), .Y(n152) );
  NAND2X1 U1042 ( .A(n239), .B(n165), .Y(n70) );
  XOR2X1 U1043 ( .A(n147), .B(n66), .Y(product_16_) );
  NAND2X1 U1044 ( .A(n235), .B(n146), .Y(n66) );
  CLKINVX1 U1045 ( .A(n145), .Y(n235) );
  XOR2X1 U1046 ( .A(n92), .B(n53), .Y(product_29_) );
  NAND2X1 U1047 ( .A(n222), .B(n91), .Y(n53) );
  CLKINVX1 U1048 ( .A(n90), .Y(n222) );
  NAND2X1 U1049 ( .A(n226), .B(n107), .Y(n57) );
  CLKINVX1 U1050 ( .A(n106), .Y(n226) );
  NAND2X1 U1051 ( .A(n228), .B(n115), .Y(n59) );
  NAND2X1 U1052 ( .A(n230), .B(n123), .Y(n61) );
  XOR2X1 U1053 ( .A(n132), .B(n63), .Y(product_19_) );
  NAND2X1 U1054 ( .A(n232), .B(n131), .Y(n63) );
  CLKINVX1 U1055 ( .A(n130), .Y(n232) );
  CLKINVX1 U1056 ( .A(n189), .Y(n188) );
  CLKINVX1 U1057 ( .A(n155), .Y(n153) );
  CLKINVX1 U1058 ( .A(n88), .Y(n86) );
  NAND2X1 U1059 ( .A(n242), .B(n184), .Y(n73) );
  XNOR2X1 U1060 ( .A(n97), .B(n54), .Y(product_28_) );
  NAND2X1 U1061 ( .A(n848), .B(n96), .Y(n54) );
  CMPR42X1 U1062 ( .A(n334), .B(n338), .C(n335), .D(n325), .ICI(n331), .S(n322), .ICO(n320), .CO(n321) );
  NOR2X1 U1063 ( .A(n183), .B(n186), .Y(n181) );
  NAND2X1 U1064 ( .A(n842), .B(n839), .Y(n190) );
  AOI21X1 U1065 ( .A0(n842), .A1(n198), .B0(n193), .Y(n191) );
  AOI21X1 U1066 ( .A0(n207), .A1(n845), .B0(n204), .Y(n202) );
  CLKINVX1 U1067 ( .A(n206), .Y(n204) );
  NOR2X2 U1068 ( .A(n375), .B(n384), .Y(n161) );
  CLKINVX1 U1069 ( .A(n96), .Y(n94) );
  AOI21X1 U1070 ( .A0(n215), .A1(n844), .B0(n212), .Y(n210) );
  CLKINVX1 U1071 ( .A(n214), .Y(n212) );
  OAI21X1 U1072 ( .A0(n216), .A1(n219), .B0(n217), .Y(n215) );
  CLKBUFX3 U1073 ( .A(b_16_), .Y(n721) );
  NAND2X1 U1074 ( .A(n857), .B(n83), .Y(n51) );
  NAND2X1 U1075 ( .A(n441), .B(n251), .Y(n83) );
  NAND2X1 U1076 ( .A(n366), .B(n374), .Y(n156) );
  NAND2X1 U1077 ( .A(n344), .B(n354), .Y(n146) );
  NAND2X1 U1078 ( .A(n312), .B(n303), .Y(n128) );
  NAND2X1 U1079 ( .A(n401), .B(n406), .Y(n178) );
  NAND2X1 U1080 ( .A(n393), .B(n400), .Y(n173) );
  NAND2X1 U1081 ( .A(n322), .B(n332), .Y(n136) );
  NAND2X1 U1082 ( .A(n407), .B(n413), .Y(n184) );
  NAND2X1 U1083 ( .A(n375), .B(n384), .Y(n162) );
  NAND2X1 U1084 ( .A(n333), .B(n343), .Y(n143) );
  NAND2X1 U1085 ( .A(n355), .B(n365), .Y(n151) );
  NAND2X1 U1086 ( .A(n313), .B(n321), .Y(n131) );
  CLKINVX1 U1087 ( .A(n208), .Y(n247) );
  XOR2X1 U1088 ( .A(n196), .B(n75), .Y(product_7_) );
  AOI21X1 U1089 ( .A0(n201), .A1(n839), .B0(n198), .Y(n196) );
  CLKINVX1 U1090 ( .A(n186), .Y(n243) );
  NAND2X1 U1091 ( .A(n224), .B(n99), .Y(n55) );
  CLKINVX1 U1092 ( .A(n98), .Y(n224) );
  XOR2X1 U1093 ( .A(n80), .B(n219), .Y(product_2_) );
  CLKINVX1 U1094 ( .A(n329), .Y(n330) );
  XNOR2X1 U1095 ( .A(n201), .B(n76), .Y(product_6_) );
  NAND2X1 U1096 ( .A(n839), .B(n200), .Y(n76) );
  CLKINVX1 U1097 ( .A(n195), .Y(n193) );
  NAND2X1 U1098 ( .A(n294), .B(n287), .Y(n120) );
  NAND2X1 U1099 ( .A(n268), .B(n264), .Y(n104) );
  NAND2X1 U1100 ( .A(n274), .B(n280), .Y(n112) );
  NAND2X1 U1101 ( .A(n302), .B(n295), .Y(n123) );
  NAND2X1 U1102 ( .A(n281), .B(n286), .Y(n115) );
  NAND2X1 U1103 ( .A(n269), .B(n273), .Y(n107) );
  NAND2X1 U1104 ( .A(n253), .B(n252), .Y(n88) );
  CLKINVX1 U1105 ( .A(n251), .Y(n252) );
  NAND2X1 U1106 ( .A(n254), .B(n255), .Y(n91) );
  OR2X1 U1107 ( .A(n441), .B(n251), .Y(n857) );
  OAI22XL U1108 ( .A0(n41), .A1(n604), .B0(n603), .B1(n755), .Y(n309) );
  OAI22XL U1109 ( .A0(n710), .A1(n4), .B0(n5), .B1(n711), .Y(n568) );
  OAI22XL U1110 ( .A0(n662), .A1(n21), .B0(n663), .B1(n24), .Y(n520) );
  CMPR42X1 U1111 ( .A(n553), .B(n420), .C(n537), .D(n416), .ICI(n417), .S(n414), .ICO(n412), .CO(n413) );
  OAI22XL U1112 ( .A0(n680), .A1(n17), .B0(n679), .B1(n759), .Y(n537) );
  CMPR42X1 U1113 ( .A(n532), .B(n380), .C(n387), .D(n378), .ICI(n383), .S(n375), .ICO(n373), .CO(n374) );
  OAI22XL U1114 ( .A0(n674), .A1(n16), .B0(n17), .B1(n675), .Y(n532) );
  OAI22XL U1115 ( .A0(n661), .A1(n24), .B0(n660), .B1(n21), .Y(n518) );
  OAI22XL U1116 ( .A0(n692), .A1(n760), .B0(n752), .B1(n693), .Y(n550) );
  CMPR42X1 U1117 ( .A(n390), .B(n549), .C(n395), .D(n391), .ICI(n388), .S(n385), .ICO(n383), .CO(n384) );
  OAI22XL U1118 ( .A0(n692), .A1(n752), .B0(n691), .B1(n760), .Y(n549) );
  CMPR42X1 U1119 ( .A(n371), .B(n361), .C(n368), .D(n358), .ICI(n364), .S(n355), .ICO(n353), .CO(n354) );
  CMPR42X1 U1120 ( .A(n379), .B(n372), .C(n377), .D(n369), .ICI(n373), .S(n366), .ICO(n364), .CO(n365) );
  CMPR42X1 U1121 ( .A(n339), .B(n560), .C(n346), .D(n342), .ICI(n336), .S(n333), .ICO(n331), .CO(n332) );
  AO21X1 U1122 ( .A0(n5), .A1(n4), .B0(n703), .Y(n560) );
  CMPR42X1 U1123 ( .A(n323), .B(n542), .C(n324), .D(n316), .ICI(n320), .S(n313), .ICO(n311), .CO(n312) );
  AO21X1 U1124 ( .A0(n752), .A1(n760), .B0(n685), .Y(n542) );
  CMPR42X1 U1125 ( .A(n314), .B(n525), .C(n306), .D(n315), .ICI(n311), .S(n303), .ICO(n301), .CO(n302) );
  OAI22XL U1126 ( .A0(n667), .A1(n16), .B0(n17), .B1(n668), .Y(n525) );
  OAI22XL U1127 ( .A0(n752), .A1(n687), .B0(n686), .B1(n760), .Y(n544) );
  OAI22XL U1128 ( .A0(n24), .A1(n658), .B0(n657), .B1(n21), .Y(n515) );
  OAI22XL U1129 ( .A0(n608), .A1(n40), .B0(n609), .B1(n41), .Y(n468) );
  OAI22XL U1130 ( .A0(n626), .A1(n748), .B0(n625), .B1(n33), .Y(n483) );
  OAI22XL U1131 ( .A0(n692), .A1(n752), .B0(n695), .B1(n760), .Y(n555) );
  OAI22XL U1132 ( .A0(n692), .A1(n760), .B0(n695), .B1(n752), .Y(n556) );
  NAND2X1 U1133 ( .A(n414), .B(n418), .Y(n187) );
  CMPR42X1 U1134 ( .A(n512), .B(n351), .C(n341), .D(n480), .ICI(n348), .S(n339), .ICO(n337), .CO(n338) );
  OAI22XL U1135 ( .A0(n654), .A1(n22), .B0(n24), .B1(n655), .Y(n512) );
  OAI22XL U1136 ( .A0(n623), .A1(n748), .B0(n622), .B1(n33), .Y(n480) );
  XNOR2X1 U1137 ( .A(n544), .B(n528), .Y(n341) );
  NAND2X1 U1138 ( .A(n419), .B(n423), .Y(n195) );
  CMPR42X1 U1139 ( .A(n317), .B(n308), .C(n449), .D(n478), .ICI(n318), .S(n306), .ICO(n304), .CO(n305) );
  OAI22XL U1140 ( .A0(n588), .A1(n48), .B0(n587), .B1(n46), .Y(n449) );
  OAI22XL U1141 ( .A0(n620), .A1(n36), .B0(n619), .B1(n34), .Y(n478) );
  NAND2X1 U1142 ( .A(n424), .B(n425), .Y(n200) );
  NAND2X1 U1143 ( .A(n575), .B(n559), .Y(n217) );
  CMPR42X1 U1144 ( .A(n481), .B(n513), .C(n467), .D(n356), .ICI(n360), .S(n347), .ICO(n345), .CO(n346) );
  OAI22XL U1145 ( .A0(n627), .A1(n748), .B0(n623), .B1(n33), .Y(n481) );
  OAI22XL U1146 ( .A0(n608), .A1(n41), .B0(n607), .B1(n755), .Y(n467) );
  OAI22XL U1147 ( .A0(n656), .A1(n24), .B0(n655), .B1(n22), .Y(n513) );
  NAND2X1 U1148 ( .A(n426), .B(n429), .Y(n206) );
  CMPR42X1 U1149 ( .A(n433), .B(n482), .C(n468), .D(n514), .ICI(n367), .S(n358), .ICO(n356), .CO(n357) );
  OAI22XL U1150 ( .A0(n625), .A1(n748), .B0(n627), .B1(n33), .Y(n482) );
  OAI22XL U1151 ( .A0(n594), .A1(n46), .B0(n48), .B1(n762), .Y(n433) );
  OAI22XL U1152 ( .A0(n656), .A1(n22), .B0(n750), .B1(n657), .Y(n514) );
  CMPR42X1 U1153 ( .A(n527), .B(n511), .C(n330), .D(n340), .ICI(n465), .S(n328), .ICO(n326), .CO(n327) );
  OAI22XL U1154 ( .A0(n606), .A1(n41), .B0(n605), .B1(n755), .Y(n465) );
  OAI22XL U1155 ( .A0(n654), .A1(n24), .B0(n653), .B1(n22), .Y(n511) );
  OR2X1 U1156 ( .A(n544), .B(n528), .Y(n340) );
  CMPR42X1 U1157 ( .A(n337), .B(n451), .C(n495), .D(n328), .ICI(n543), .S(n325), .ICO(n323), .CO(n324) );
  OAI22XL U1158 ( .A0(n685), .A1(n760), .B0(n752), .B1(n686), .Y(n543) );
  OAI22XL U1159 ( .A0(n638), .A1(n29), .B0(n637), .B1(n28), .Y(n495) );
  OAI22XL U1160 ( .A0(n590), .A1(n48), .B0(n589), .B1(n46), .Y(n451) );
  CMPR42X1 U1161 ( .A(n326), .B(n464), .C(n479), .D(n327), .ICI(n319), .S(n316), .ICO(n314), .CO(n315) );
  OAI22XL U1162 ( .A0(n605), .A1(n41), .B0(n604), .B1(n755), .Y(n464) );
  OAI22XL U1163 ( .A0(n620), .A1(n34), .B0(n748), .B1(n621), .Y(n479) );
  CMPR42X1 U1164 ( .A(n350), .B(n561), .C(n357), .D(n353), .ICI(n347), .S(n344), .ICO(n342), .CO(n343) );
  OAI22XL U1165 ( .A0(n703), .A1(n4), .B0(n5), .B1(n704), .Y(n561) );
  CMPR42X1 U1166 ( .A(n567), .B(n519), .C(n408), .D(n405), .ICI(n404), .S(n401), .ICO(n399), .CO(n400) );
  OAI22XL U1167 ( .A0(n662), .A1(n24), .B0(n661), .B1(n21), .Y(n519) );
  OAI22XL U1168 ( .A0(n710), .A1(n753), .B0(n709), .B1(n4), .Y(n567) );
  NAND2X1 U1169 ( .A(n430), .B(n431), .Y(n209) );
  CMPR42X1 U1170 ( .A(n510), .B(n329), .C(n526), .D(n494), .ICI(n450), .S(n319), .ICO(n317), .CO(n318) );
  OAI22XL U1171 ( .A0(n636), .A1(n28), .B0(n29), .B1(n637), .Y(n494) );
  OAI22XL U1172 ( .A0(n17), .A1(n669), .B0(n668), .B1(n16), .Y(n526) );
  OAI22XL U1173 ( .A0(n589), .A1(n48), .B0(n588), .B1(n46), .Y(n450) );
  CMPR42X1 U1174 ( .A(n466), .B(n496), .C(n452), .D(n349), .ICI(n345), .S(n336), .ICO(n334), .CO(n335) );
  OAI22XL U1175 ( .A0(n607), .A1(n41), .B0(n606), .B1(n755), .Y(n466) );
  OAI22XL U1176 ( .A0(n590), .A1(n46), .B0(n591), .B1(n48), .Y(n452) );
  OAI22XL U1177 ( .A0(n638), .A1(n28), .B0(n29), .B1(n639), .Y(n496) );
  OAI22XL U1178 ( .A0(n708), .A1(n4), .B0(n753), .B1(n709), .Y(n566) );
  ADDFXL U1179 ( .A(n533), .B(n565), .CI(n471), .CO(n389), .S(n390) );
  OAI22XL U1180 ( .A0(n708), .A1(n5), .B0(n707), .B1(n4), .Y(n565) );
  NOR2BX1 U1181 ( .AN(n49), .B(n40), .Y(n471) );
  CLKINVX1 U1182 ( .A(n81), .Y(product_1_) );
  OAI22XL U1183 ( .A0(n586), .A1(n48), .B0(n46), .B1(n585), .Y(n291) );
  CMPR42X1 U1184 ( .A(n276), .B(n446), .C(n283), .D(n489), .ICI(n279), .S(n274), .ICO(n272), .CO(n273) );
  OAI22XL U1185 ( .A0(n584), .A1(n48), .B0(n46), .B1(n583), .Y(n446) );
  OAI22XL U1186 ( .A0(n631), .A1(n28), .B0(n749), .B1(n632), .Y(n489) );
  CMPR42X1 U1187 ( .A(n447), .B(n284), .C(n289), .D(n506), .ICI(n285), .S(n281), .ICO(n279), .CO(n280) );
  OAI22XL U1188 ( .A0(n584), .A1(n46), .B0(n48), .B1(n585), .Y(n447) );
  AO21X1 U1189 ( .A0(n24), .A1(n22), .B0(n649), .Y(n506) );
  CMPR42X1 U1190 ( .A(n445), .B(n271), .C(n275), .D(n272), .ICI(n488), .S(n269), .ICO(n267), .CO(n268) );
  OAI22XL U1191 ( .A0(n582), .A1(n46), .B0(n48), .B1(n583), .Y(n445) );
  CMPR42X1 U1192 ( .A(n462), .B(n290), .C(n507), .D(n297), .ICI(n293), .S(n287), .ICO(n285), .CO(n286) );
  OAI22XL U1193 ( .A0(n602), .A1(n42), .B0(n601), .B1(n40), .Y(n462) );
  OAI22XL U1194 ( .A0(n649), .A1(n22), .B0(n24), .B1(n650), .Y(n507) );
  CMPR42X1 U1195 ( .A(n304), .B(n524), .C(n298), .D(n305), .ICI(n301), .S(n295), .ICO(n293), .CO(n294) );
  AO21X1 U1196 ( .A0(n17), .A1(n16), .B0(n667), .Y(n524) );
  CMPR42X1 U1197 ( .A(n444), .B(n266), .C(n270), .D(n267), .ICI(n473), .S(n264), .ICO(n262), .CO(n263) );
  OAI22XL U1198 ( .A0(n582), .A1(n48), .B0(n46), .B1(n581), .Y(n444) );
  CLKINVX1 U1199 ( .A(n265), .Y(n266) );
  OAI22XL U1200 ( .A0(n613), .A1(n34), .B0(n36), .B1(n614), .Y(n473) );
  CLKBUFX3 U1201 ( .A(b_15_), .Y(n722) );
  CMPR42X1 U1202 ( .A(n477), .B(n300), .C(n307), .D(n448), .ICI(n463), .S(n298), .ICO(n296), .CO(n297) );
  OAI22XL U1203 ( .A0(n618), .A1(n34), .B0(n36), .B1(n619), .Y(n477) );
  OAI22XL U1204 ( .A0(n602), .A1(n40), .B0(n41), .B1(n603), .Y(n463) );
  OAI22XL U1205 ( .A0(n587), .A1(n48), .B0(n586), .B1(n46), .Y(n448) );
  ADDFXL U1206 ( .A(n460), .B(n278), .CI(n282), .CO(n275), .S(n276) );
  OAI22XL U1207 ( .A0(n600), .A1(n42), .B0(n599), .B1(n40), .Y(n460) );
  CLKINVX1 U1208 ( .A(n277), .Y(n278) );
  CLKINVX1 U1209 ( .A(n43), .Y(n762) );
  XNOR2X1 U1210 ( .A(n721), .B(n43), .Y(n577) );
  CLKINVX1 U1211 ( .A(n257), .Y(n258) );
  OAI22XL U1212 ( .A0(n595), .A1(n40), .B0(n42), .B1(n596), .Y(n457) );
  OAI22XL U1213 ( .A0(n579), .A1(n48), .B0(n46), .B1(n578), .Y(n442) );
  NAND2X1 U1214 ( .A(n256), .B(n260), .Y(n96) );
  NAND2X1 U1215 ( .A(n261), .B(n263), .Y(n99) );
  XNOR2X1 U1216 ( .A(n43), .B(n722), .Y(n578) );
  OAI22X1 U1217 ( .A0(n717), .A1(n4), .B0(n5), .B1(n718), .Y(n575) );
  OAI22X1 U1218 ( .A0(n719), .A1(n5), .B0(n718), .B1(n4), .Y(n576) );
  XNOR2X1 U1219 ( .A(n49), .B(n1), .Y(n719) );
  CMPR42X1 U1220 ( .A(n553), .B(n522), .C(n421), .D(n538), .ICI(n422), .S(n419), .ICO(n417), .CO(n418) );
  OAI22XL U1221 ( .A0(n680), .A1(n16), .B0(n681), .B1(n17), .Y(n538) );
  NOR2BX1 U1222 ( .AN(n49), .B(n21), .Y(n523) );
  XNOR2X1 U1223 ( .A(n1), .B(b_12_), .Y(n707) );
  XNOR2X1 U1224 ( .A(n1), .B(b_10_), .Y(n709) );
  XNOR2X1 U1225 ( .A(n7), .B(n722), .Y(n691) );
  XNOR2X1 U1226 ( .A(n1), .B(n722), .Y(n704) );
  XNOR2X1 U1227 ( .A(n1), .B(n729), .Y(n711) );
  XNOR2X1 U1228 ( .A(n734), .B(n1), .Y(n716) );
  XNOR2X1 U1229 ( .A(b_11_), .B(n1), .Y(n708) );
  XNOR2X1 U1230 ( .A(n728), .B(n1), .Y(n710) );
  XNOR2X1 U1231 ( .A(b_11_), .B(n7), .Y(n690) );
  XNOR2X1 U1232 ( .A(n733), .B(n13), .Y(n679) );
  XNOR2X1 U1233 ( .A(n735), .B(n19), .Y(n663) );
  XNOR2X1 U1234 ( .A(b_5_), .B(n13), .Y(n678) );
  XNOR2X1 U1235 ( .A(b_7_), .B(n7), .Y(n694) );
  XNOR2X1 U1236 ( .A(n723), .B(n1), .Y(n705) );
  XNOR2X1 U1237 ( .A(b_7_), .B(n31), .Y(n622) );
  XNOR2X1 U1238 ( .A(n721), .B(n1), .Y(n703) );
  CLKINVX1 U1239 ( .A(n7), .Y(n768) );
  OAI22XL U1240 ( .A0(n17), .A1(n670), .B0(n669), .B1(n16), .Y(n527) );
  ADDHXL U1241 ( .A(n564), .B(n548), .CO(n381), .S(n382) );
  OAI22XL U1242 ( .A0(n753), .A1(n707), .B0(n706), .B1(n4), .Y(n564) );
  OAI22XL U1243 ( .A0(n690), .A1(n760), .B0(n752), .B1(n691), .Y(n548) );
  ADDHXL U1244 ( .A(n546), .B(n562), .CO(n362), .S(n363) );
  OAI22XL U1245 ( .A0(n5), .A1(n705), .B0(n704), .B1(n4), .Y(n562) );
  OAI22XL U1246 ( .A0(n752), .A1(n689), .B0(n688), .B1(n760), .Y(n546) );
  ADDHXL U1247 ( .A(n497), .B(n545), .CO(n351), .S(n352) );
  OAI22XL U1248 ( .A0(n752), .A1(n688), .B0(n687), .B1(n760), .Y(n545) );
  OAI22XL U1249 ( .A0(n29), .A1(n640), .B0(n639), .B1(n28), .Y(n497) );
  CLKINVX1 U1250 ( .A(n25), .Y(n765) );
  CLKINVX1 U1251 ( .A(n13), .Y(n767) );
  CMPR42X1 U1252 ( .A(n530), .B(n363), .C(n370), .D(n498), .ICI(n454), .S(n361), .ICO(n359), .CO(n360) );
  OAI22XL U1253 ( .A0(n593), .A1(n48), .B0(n46), .B1(n592), .Y(n454) );
  OAI22XL U1254 ( .A0(n672), .A1(n16), .B0(n17), .B1(n673), .Y(n530) );
  OAI22XL U1255 ( .A0(n641), .A1(n29), .B0(n640), .B1(n28), .Y(n498) );
  CMPR42X1 U1256 ( .A(n515), .B(n563), .C(n547), .D(n381), .ICI(n499), .S(n372), .ICO(n370), .CO(n371) );
  OAI22XL U1257 ( .A0(n642), .A1(n29), .B0(n641), .B1(n28), .Y(n499) );
  OAI22XL U1258 ( .A0(n753), .A1(n706), .B0(n705), .B1(n4), .Y(n563) );
  OAI22XL U1259 ( .A0(n690), .A1(n752), .B0(n689), .B1(n760), .Y(n547) );
  OAI22XL U1260 ( .A0(n644), .A1(n28), .B0(n645), .B1(n29), .Y(n502) );
  CMPR42X1 U1261 ( .A(n551), .B(n487), .C(n503), .D(n535), .ICI(n410), .S(n404), .ICO(n402), .CO(n403) );
  OAI22XL U1262 ( .A0(n678), .A1(n17), .B0(n678), .B1(n16), .Y(n535) );
  OAI22XL U1263 ( .A0(n645), .A1(n28), .B0(n29), .B1(n646), .Y(n503) );
  CMPR42X1 U1264 ( .A(n485), .B(n517), .C(n397), .D(n501), .ICI(n394), .S(n388), .ICO(n386), .CO(n387) );
  OAI22XL U1265 ( .A0(n644), .A1(n29), .B0(n643), .B1(n28), .Y(n501) );
  OAI22XL U1266 ( .A0(n627), .A1(n33), .B0(n748), .B1(n628), .Y(n485) );
  OAI22XL U1267 ( .A0(n626), .A1(n33), .B0(n627), .B1(n748), .Y(n484) );
  CMPR42X1 U1268 ( .A(n455), .B(n469), .C(n483), .D(n531), .ICI(n376), .S(n369), .ICO(n367), .CO(n368) );
  NOR2BX1 U1269 ( .AN(n49), .B(n46), .Y(n455) );
  OAI22XL U1270 ( .A0(n609), .A1(n40), .B0(n41), .B1(n610), .Y(n469) );
  OAI22XL U1271 ( .A0(n674), .A1(n17), .B0(n673), .B1(n16), .Y(n531) );
  CMPR42X1 U1272 ( .A(n529), .B(n352), .C(n362), .D(n453), .ICI(n359), .S(n350), .ICO(n348), .CO(n349) );
  OAI22XL U1273 ( .A0(n672), .A1(n17), .B0(n671), .B1(n16), .Y(n529) );
  OAI22XL U1274 ( .A0(n591), .A1(n46), .B0(n48), .B1(n592), .Y(n453) );
  CLKBUFX3 U1275 ( .A(n754), .Y(n46) );
  CLKBUFX3 U1276 ( .A(n759), .Y(n16) );
  CLKBUFX3 U1277 ( .A(n756), .Y(n34) );
  CLKBUFX3 U1278 ( .A(n756), .Y(n33) );
  CLKBUFX3 U1279 ( .A(n761), .Y(n4) );
  ADDFXL U1280 ( .A(n509), .B(n493), .CI(n310), .CO(n307), .S(n308) );
  OAI22XL U1281 ( .A0(n24), .A1(n652), .B0(n651), .B1(n22), .Y(n509) );
  OAI22XL U1282 ( .A0(n636), .A1(n29), .B0(n635), .B1(n28), .Y(n493) );
  CLKINVX1 U1283 ( .A(n309), .Y(n310) );
  OAI22XL U1284 ( .A0(n612), .A1(n40), .B0(n42), .B1(n763), .Y(n434) );
  CLKINVX1 U1285 ( .A(n37), .Y(n763) );
  CLKBUFX3 U1286 ( .A(n747), .Y(n41) );
  CLKBUFX3 U1287 ( .A(n748), .Y(n36) );
  ADDFXL U1288 ( .A(n569), .B(n505), .CI(n521), .CO(n415), .S(n416) );
  OAI22XL U1289 ( .A0(n5), .A1(n712), .B0(n711), .B1(n4), .Y(n569) );
  NOR2BX1 U1290 ( .AN(n49), .B(n28), .Y(n505) );
  OAI22XL U1291 ( .A0(n647), .A1(n29), .B0(n646), .B1(n28), .Y(n504) );
  CLKINVX1 U1292 ( .A(n31), .Y(n764) );
  OAI22XL U1293 ( .A0(n24), .A1(n653), .B0(n652), .B1(n22), .Y(n510) );
  CMPR42X1 U1294 ( .A(n291), .B(n475), .C(n490), .D(n461), .ICI(n288), .S(n284), .ICO(n282), .CO(n283) );
  OAI22XL U1295 ( .A0(n600), .A1(n40), .B0(n42), .B1(n601), .Y(n461) );
  OAI22XL U1296 ( .A0(n749), .A1(n633), .B0(n632), .B1(n28), .Y(n490) );
  OAI22XL U1297 ( .A0(n36), .A1(n617), .B0(n616), .B1(n34), .Y(n475) );
  CMPR42X1 U1298 ( .A(n491), .B(n292), .C(n476), .D(n299), .ICI(n296), .S(n290), .ICO(n288), .CO(n289) );
  OAI22XL U1299 ( .A0(n618), .A1(n36), .B0(n617), .B1(n34), .Y(n476) );
  OAI22XL U1300 ( .A0(n29), .A1(n634), .B0(n633), .B1(n28), .Y(n491) );
  CLKINVX1 U1301 ( .A(n291), .Y(n292) );
  ADDFXL U1302 ( .A(n474), .B(n459), .CI(n277), .CO(n270), .S(n271) );
  OAI22XL U1303 ( .A0(n36), .A1(n615), .B0(n614), .B1(n34), .Y(n474) );
  OAI22XL U1304 ( .A0(n42), .A1(n599), .B0(n598), .B1(n40), .Y(n459) );
  ADDFXL U1305 ( .A(n309), .B(n492), .CI(n508), .CO(n299), .S(n300) );
  OAI22XL U1306 ( .A0(n24), .A1(n651), .B0(n650), .B1(n22), .Y(n508) );
  OAI22XL U1307 ( .A0(n29), .A1(n635), .B0(n634), .B1(n28), .Y(n492) );
  CMPR42X1 U1308 ( .A(n443), .B(n458), .C(n265), .D(n262), .ICI(n472), .S(n261), .ICO(n259), .CO(n260) );
  OAI22XL U1309 ( .A0(n42), .A1(n597), .B0(n596), .B1(n40), .Y(n458) );
  OAI22XL U1310 ( .A0(n48), .A1(n581), .B0(n46), .B1(n580), .Y(n443) );
  XNOR2X2 U1311 ( .A(a_11_), .B(a_12_), .Y(n755) );
  XNOR2X1 U1312 ( .A(n1), .B(n724), .Y(n706) );
  XNOR2X1 U1313 ( .A(n1), .B(n736), .Y(n718) );
  XNOR2X1 U1314 ( .A(n13), .B(n736), .Y(n682) );
  XNOR2X1 U1315 ( .A(n31), .B(n736), .Y(n628) );
  XNOR2X1 U1316 ( .A(n25), .B(n736), .Y(n646) );
  XNOR2X1 U1317 ( .A(n37), .B(n736), .Y(n610) );
  NAND2X1 U1318 ( .A(n743), .B(n759), .Y(n751) );
  XOR2X1 U1319 ( .A(a_7_), .B(a_6_), .Y(n742) );
  XOR2X1 U1320 ( .A(a_9_), .B(a_8_), .Y(n741) );
  XOR2X1 U1321 ( .A(a_11_), .B(a_10_), .Y(n740) );
  NAND2X1 U1322 ( .A(n739), .B(n755), .Y(n747) );
  XOR2X1 U1323 ( .A(a_13_), .B(a_12_), .Y(n739) );
  XOR2X1 U1324 ( .A(a_3_), .B(a_2_), .Y(n744) );
  NAND2X1 U1325 ( .A(n754), .B(n738), .Y(n746) );
  XOR2X1 U1326 ( .A(a_14_), .B(a_15_), .Y(n738) );
  NAND2X1 U1327 ( .A(n745), .B(n761), .Y(n753) );
  XOR2X1 U1328 ( .A(a_0_), .B(a_1_), .Y(n745) );
  XNOR2X1 U1329 ( .A(n31), .B(n724), .Y(n616) );
  XNOR2X1 U1330 ( .A(n43), .B(n736), .Y(n592) );
  XNOR2X1 U1331 ( .A(n37), .B(n724), .Y(n598) );
endmodule


module FFT_ultrafast2_shift_DW01_add_22 ( A, B, SUM_31_, SUM_30_, SUM_29_, 
        SUM_28_, SUM_27_, SUM_26_, SUM_25_, SUM_24_, SUM_23_, SUM_22_, SUM_21_, 
        SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_ );
  input [31:0] A;
  input [31:0] B;
  output SUM_31_, SUM_30_, SUM_29_, SUM_28_, SUM_27_, SUM_26_, SUM_25_,
         SUM_24_, SUM_23_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_,
         SUM_17_, SUM_16_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n21, n23, n24, n25, n26, n27, n29, n31, n32, n33, n34, n35, n37,
         n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51, n53, n55, n56,
         n57, n58, n59, n61, n63, n64, n65, n66, n67, n69, n71, n72, n73, n74,
         n76, n78, n79, n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n121, n124, n125, n127, n128, n129, n132, n133, n135, n136, n137,
         n140, n141, n143, n144, n145, n148, n149, n151, n154, n156, n158,
         n160, n162, n164, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276;

  OAI21X1 U187 ( .A0(n111), .A1(n121), .B0(n112), .Y(n110) );
  AOI21X1 U188 ( .A0(n275), .A1(n267), .B0(n265), .Y(n112) );
  OR2X1 U189 ( .A(B[13]), .B(A[13]), .Y(n273) );
  NAND2X1 U190 ( .A(B[28]), .B(A[28]), .Y(n31) );
  OR2X1 U191 ( .A(B[18]), .B(A[18]), .Y(n262) );
  OR2X1 U192 ( .A(A[17]), .B(B[17]), .Y(n256) );
  NAND2X1 U193 ( .A(A[16]), .B(B[16]), .Y(n83) );
  BUFX3 U194 ( .A(A[4]), .Y(n254) );
  OR2X1 U195 ( .A(A[16]), .B(B[16]), .Y(n255) );
  OR2X1 U196 ( .A(B[30]), .B(A[30]), .Y(n257) );
  OR2X1 U197 ( .A(B[28]), .B(A[28]), .Y(n258) );
  OR2X1 U198 ( .A(B[20]), .B(A[20]), .Y(n259) );
  OR2XL U199 ( .A(B[22]), .B(A[22]), .Y(n260) );
  OR2X1 U200 ( .A(B[26]), .B(A[26]), .Y(n261) );
  OR2X1 U201 ( .A(B[24]), .B(A[24]), .Y(n263) );
  AND2X2 U202 ( .A(B[13]), .B(A[13]), .Y(n264) );
  AND2X2 U203 ( .A(B[9]), .B(A[9]), .Y(n265) );
  AND2X2 U204 ( .A(A[12]), .B(B[12]), .Y(n266) );
  AND2X2 U205 ( .A(A[8]), .B(B[8]), .Y(n267) );
  OR2X2 U206 ( .A(B[9]), .B(A[9]), .Y(n275) );
  OR2X1 U207 ( .A(A[8]), .B(B[8]), .Y(n270) );
  AOI21X1 U208 ( .A0(n273), .A1(n266), .B0(n264), .Y(n94) );
  NAND2X1 U209 ( .A(B[26]), .B(A[26]), .Y(n39) );
  NOR2XL U210 ( .A(A[10]), .B(B[10]), .Y(n108) );
  AO21X4 U211 ( .A0(n24), .A1(n257), .B0(n21), .Y(n268) );
  OAI21X2 U212 ( .A0(n43), .A1(n41), .B0(n42), .Y(n40) );
  OAI21X2 U213 ( .A0(n51), .A1(n49), .B0(n50), .Y(n48) );
  XNOR2X1 U214 ( .A(n268), .B(n1), .Y(SUM_31_) );
  NAND2XL U215 ( .A(A[7]), .B(B[7]), .Y(n125) );
  OAI21X1 U216 ( .A0(n85), .A1(n73), .B0(n74), .Y(n72) );
  AOI21X1 U217 ( .A0(n256), .A1(n81), .B0(n76), .Y(n74) );
  INVX1 U218 ( .A(n78), .Y(n76) );
  NOR2X1 U219 ( .A(n88), .B(n90), .Y(n86) );
  NAND2X1 U220 ( .A(B[30]), .B(A[30]), .Y(n23) );
  OAI21X2 U221 ( .A0(n35), .A1(n33), .B0(n34), .Y(n32) );
  OAI21X1 U222 ( .A0(n88), .A1(n91), .B0(n89), .Y(n87) );
  OAI21X1 U223 ( .A0(n103), .A1(n93), .B0(n94), .Y(n92) );
  NAND2XL U224 ( .A(A[6]), .B(B[6]), .Y(n128) );
  NAND2XL U225 ( .A(A[1]), .B(B[1]), .Y(n149) );
  OAI21X1 U226 ( .A0(n59), .A1(n57), .B0(n58), .Y(n56) );
  OAI21X1 U227 ( .A0(n67), .A1(n65), .B0(n66), .Y(n64) );
  NOR2X2 U228 ( .A(A[29]), .B(B[29]), .Y(n25) );
  NAND2X1 U229 ( .A(A[29]), .B(B[29]), .Y(n26) );
  OA21XL U230 ( .A0(n271), .A1(n132), .B0(n133), .Y(n129) );
  OA21XL U231 ( .A0(n137), .A1(n135), .B0(n136), .Y(n271) );
  NAND2X1 U232 ( .A(A[27]), .B(B[27]), .Y(n34) );
  OR2X1 U233 ( .A(A[31]), .B(B[31]), .Y(n276) );
  OAI21X2 U234 ( .A0(n27), .A1(n25), .B0(n26), .Y(n24) );
  XNOR2XL U235 ( .A(n48), .B(n8), .Y(SUM_24_) );
  NAND2XL U236 ( .A(n263), .B(n47), .Y(n8) );
  XOR2XL U237 ( .A(n67), .B(n13), .Y(SUM_19_) );
  NAND2XL U238 ( .A(n164), .B(n66), .Y(n13) );
  XNOR2XL U239 ( .A(n72), .B(n14), .Y(SUM_18_) );
  NAND2XL U240 ( .A(n262), .B(n71), .Y(n14) );
  NAND2XL U241 ( .A(n256), .B(n78), .Y(n15) );
  AOI21XL U242 ( .A0(n84), .A1(n255), .B0(n81), .Y(n79) );
  INVXL U243 ( .A(n85), .Y(n84) );
  NOR2X1 U244 ( .A(A[21]), .B(B[21]), .Y(n57) );
  NOR2X1 U245 ( .A(A[25]), .B(B[25]), .Y(n41) );
  NOR2X1 U246 ( .A(A[23]), .B(B[23]), .Y(n49) );
  NOR2X1 U247 ( .A(A[19]), .B(B[19]), .Y(n65) );
  NAND2XL U248 ( .A(A[15]), .B(B[15]), .Y(n89) );
  OR2X1 U249 ( .A(A[12]), .B(B[12]), .Y(n269) );
  NOR2X1 U250 ( .A(A[27]), .B(B[27]), .Y(n33) );
  NAND2XL U251 ( .A(A[11]), .B(B[11]), .Y(n107) );
  NAND2XL U252 ( .A(B[2]), .B(A[2]), .Y(n144) );
  XNOR2X1 U253 ( .A(n24), .B(n2), .Y(SUM_30_) );
  NAND2X1 U254 ( .A(n257), .B(n23), .Y(n2) );
  XNOR2X1 U255 ( .A(n40), .B(n6), .Y(SUM_26_) );
  NAND2X1 U256 ( .A(n261), .B(n39), .Y(n6) );
  AOI21X1 U257 ( .A0(n72), .A1(n262), .B0(n69), .Y(n67) );
  CLKINVX1 U258 ( .A(n71), .Y(n69) );
  AOI21X1 U259 ( .A0(n64), .A1(n259), .B0(n61), .Y(n59) );
  CLKINVX1 U260 ( .A(n63), .Y(n61) );
  AOI21X1 U261 ( .A0(n56), .A1(n260), .B0(n53), .Y(n51) );
  CLKINVX1 U262 ( .A(n55), .Y(n53) );
  AOI21X1 U263 ( .A0(n48), .A1(n263), .B0(n45), .Y(n43) );
  CLKINVX1 U264 ( .A(n47), .Y(n45) );
  AOI21X1 U265 ( .A0(n40), .A1(n261), .B0(n37), .Y(n35) );
  CLKINVX1 U266 ( .A(n39), .Y(n37) );
  NAND2X1 U267 ( .A(n255), .B(n256), .Y(n73) );
  XOR2X1 U268 ( .A(n27), .B(n3), .Y(SUM_29_) );
  NAND2X1 U269 ( .A(n154), .B(n26), .Y(n3) );
  CLKINVX1 U270 ( .A(n25), .Y(n154) );
  XOR2X1 U271 ( .A(n43), .B(n7), .Y(SUM_25_) );
  NAND2X1 U272 ( .A(n158), .B(n42), .Y(n7) );
  CLKINVX1 U273 ( .A(n41), .Y(n158) );
  CLKINVX1 U274 ( .A(n83), .Y(n81) );
  CLKINVX1 U275 ( .A(n23), .Y(n21) );
  XNOR2X1 U276 ( .A(n56), .B(n10), .Y(SUM_22_) );
  NAND2X1 U277 ( .A(n260), .B(n55), .Y(n10) );
  XNOR2X1 U278 ( .A(n64), .B(n12), .Y(SUM_20_) );
  NAND2X1 U279 ( .A(n259), .B(n63), .Y(n12) );
  XOR2X1 U280 ( .A(n51), .B(n9), .Y(SUM_23_) );
  NAND2X1 U281 ( .A(n160), .B(n50), .Y(n9) );
  CLKINVX1 U282 ( .A(n49), .Y(n160) );
  XOR2X1 U283 ( .A(n59), .B(n11), .Y(SUM_21_) );
  NAND2X1 U284 ( .A(n162), .B(n58), .Y(n11) );
  CLKINVX1 U285 ( .A(n57), .Y(n162) );
  CLKINVX1 U286 ( .A(n65), .Y(n164) );
  XOR2X1 U287 ( .A(n79), .B(n15), .Y(SUM_17_) );
  XNOR2X1 U288 ( .A(n84), .B(n16), .Y(SUM_16_) );
  NAND2X1 U289 ( .A(n255), .B(n83), .Y(n16) );
  AOI21X1 U290 ( .A0(n92), .A1(n86), .B0(n87), .Y(n85) );
  XNOR2X1 U291 ( .A(n32), .B(n4), .Y(SUM_28_) );
  NAND2X1 U292 ( .A(n258), .B(n31), .Y(n4) );
  AOI21X1 U293 ( .A0(n32), .A1(n258), .B0(n29), .Y(n27) );
  CLKINVX1 U294 ( .A(n31), .Y(n29) );
  AOI21X1 U295 ( .A0(n104), .A1(n110), .B0(n105), .Y(n103) );
  NOR2X1 U296 ( .A(n106), .B(n108), .Y(n104) );
  OAI21XL U297 ( .A0(n106), .A1(n109), .B0(n107), .Y(n105) );
  OA21XL U298 ( .A0(n272), .A1(n124), .B0(n125), .Y(n121) );
  OA21XL U299 ( .A0(n129), .A1(n127), .B0(n128), .Y(n272) );
  NOR2X1 U300 ( .A(A[15]), .B(B[15]), .Y(n88) );
  XOR2X1 U301 ( .A(n35), .B(n5), .Y(SUM_27_) );
  NAND2X1 U302 ( .A(n156), .B(n34), .Y(n5) );
  CLKINVX1 U303 ( .A(n33), .Y(n156) );
  NAND2X1 U304 ( .A(A[17]), .B(B[17]), .Y(n78) );
  NAND2X1 U305 ( .A(B[24]), .B(A[24]), .Y(n47) );
  NAND2X1 U306 ( .A(B[22]), .B(A[22]), .Y(n55) );
  NAND2X1 U307 ( .A(B[20]), .B(A[20]), .Y(n63) );
  NAND2X1 U308 ( .A(B[18]), .B(A[18]), .Y(n71) );
  NAND2X1 U309 ( .A(A[25]), .B(B[25]), .Y(n42) );
  NAND2X1 U310 ( .A(A[23]), .B(B[23]), .Y(n50) );
  NAND2X1 U311 ( .A(A[21]), .B(B[21]), .Y(n58) );
  NAND2X1 U312 ( .A(A[19]), .B(B[19]), .Y(n66) );
  NOR2X1 U313 ( .A(B[14]), .B(A[14]), .Y(n90) );
  NAND2X1 U314 ( .A(n276), .B(n18), .Y(n1) );
  NAND2X1 U315 ( .A(B[14]), .B(A[14]), .Y(n91) );
  OA21XL U316 ( .A0(n274), .A1(n140), .B0(n141), .Y(n137) );
  OA21XL U317 ( .A0(n145), .A1(n143), .B0(n144), .Y(n274) );
  NOR2X1 U318 ( .A(A[11]), .B(B[11]), .Y(n106) );
  NOR2X1 U319 ( .A(A[3]), .B(B[3]), .Y(n140) );
  NOR2X1 U320 ( .A(B[5]), .B(A[5]), .Y(n132) );
  NOR2X1 U321 ( .A(A[7]), .B(B[7]), .Y(n124) );
  NAND2X1 U322 ( .A(A[3]), .B(B[3]), .Y(n141) );
  NOR2X1 U323 ( .A(B[2]), .B(A[2]), .Y(n143) );
  NOR2X1 U324 ( .A(A[6]), .B(B[6]), .Y(n127) );
  NOR2X1 U325 ( .A(n254), .B(B[4]), .Y(n135) );
  NAND2X1 U326 ( .A(A[10]), .B(B[10]), .Y(n109) );
  NAND2X1 U327 ( .A(A[31]), .B(B[31]), .Y(n18) );
  NAND2X1 U328 ( .A(B[5]), .B(A[5]), .Y(n133) );
  NAND2X1 U329 ( .A(n254), .B(B[4]), .Y(n136) );
  NAND2X1 U330 ( .A(n275), .B(n270), .Y(n111) );
  NAND2X1 U331 ( .A(n273), .B(n269), .Y(n93) );
  OA21XL U332 ( .A0(n148), .A1(n151), .B0(n149), .Y(n145) );
  NOR2X1 U333 ( .A(A[1]), .B(B[1]), .Y(n148) );
  NAND2X1 U334 ( .A(A[0]), .B(B[0]), .Y(n151) );
endmodule


module FFT_ultrafast2_shift_DW_mult_uns_11 ( a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_8_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, a_0_, 
        b_16_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_, 
        b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_, product_31_, product_30_, 
        product_29_, product_28_, product_27_, product_26_, product_25_, 
        product_24_, product_23_, product_22_, product_21_, product_20_, 
        product_19_, product_18_, product_17_, product_16_, product_15_, 
        product_14_, product_13_, product_12_, product_11_, product_10_, 
        product_9_, product_8_, product_7_, product_6_, product_5_, product_4_, 
        product_3_, product_2_, product_1_, product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_8_, a_7_, a_6_, a_5_,
         a_4_, a_3_, a_2_, a_1_, a_0_, b_16_, b_15_, b_14_, b_13_, b_12_,
         b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_,
         b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_1_, product_0_;
  wire   n1, n3, n5, n7, n9, n10, n11, n12, n13, n15, n16, n17, n19, n21, n22,
         n24, n25, n27, n28, n29, n31, n33, n34, n35, n36, n37, n40, n42, n43,
         n46, n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n83, n86, n88, n89, n90, n91, n92, n94,
         n96, n97, n98, n99, n100, n102, n104, n105, n106, n107, n108, n110,
         n112, n113, n114, n115, n116, n118, n120, n121, n122, n123, n124,
         n126, n128, n129, n130, n131, n132, n134, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n171, n173, n174,
         n176, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n193, n195, n196, n198, n200, n201, n202,
         n204, n206, n207, n208, n209, n210, n212, n214, n215, n216, n217,
         n218, n219, n222, n224, n226, n228, n230, n232, n234, n235, n236,
         n238, n239, n242, n243, n247, n249, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n728, n729, n730, n731,
         n732, n733, n735, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859;

  XNOR2X1 U699 ( .A(n735), .B(n7), .Y(n699) );
  CLKBUFX4 U700 ( .A(b_2_), .Y(n735) );
  OAI21X1 U701 ( .A0(n92), .A1(n90), .B0(n91), .Y(n89) );
  AOI21X2 U702 ( .A0(n97), .A1(n850), .B0(n94), .Y(n92) );
  OAI21X1 U703 ( .A0(n166), .A1(n164), .B0(n165), .Y(n163) );
  INVXL U704 ( .A(n167), .Y(n166) );
  XNOR2X2 U705 ( .A(n185), .B(n73), .Y(product_9_) );
  OAI21X1 U706 ( .A0(n188), .A1(n186), .B0(n187), .Y(n185) );
  BUFX12 U707 ( .A(n751), .Y(n17) );
  OAI22X1 U708 ( .A0(n697), .A1(n11), .B0(n696), .B1(n9), .Y(n554) );
  BUFX6 U709 ( .A(n576), .Y(n838) );
  OAI22X1 U710 ( .A0(n719), .A1(n5), .B0(n718), .B1(n3), .Y(n576) );
  ADDFX2 U711 ( .A(n536), .B(n504), .CI(n411), .CO(n408), .S(n409) );
  ADDHX1 U712 ( .A(n552), .B(n436), .CO(n410), .S(n411) );
  OAI21X4 U713 ( .A0(n116), .A1(n114), .B0(n115), .Y(n113) );
  AOI21X4 U714 ( .A0(n121), .A1(n847), .B0(n118), .Y(n116) );
  NAND2X2 U715 ( .A(n838), .B(n440), .Y(n219) );
  OAI22X1 U716 ( .A0(n720), .A1(n3), .B0(n5), .B1(n769), .Y(n440) );
  OAI22XL U717 ( .A0(n716), .A1(n3), .B0(n717), .B1(n5), .Y(n574) );
  CMPR42X1 U718 ( .A(n415), .B(n520), .C(n568), .D(n409), .ICI(n412), .S(n407), 
        .ICO(n405), .CO(n406) );
  NOR2X2 U719 ( .A(n407), .B(n413), .Y(n183) );
  OAI21X1 U720 ( .A0(n190), .A1(n202), .B0(n191), .Y(n189) );
  CMPR42X1 U721 ( .A(n554), .B(n522), .C(n421), .D(n538), .ICI(n422), .S(n419), 
        .ICO(n417), .CO(n418) );
  OAI22XL U722 ( .A0(n17), .A1(n676), .B0(n675), .B1(n15), .Y(n533) );
  XNOR2X1 U723 ( .A(n7), .B(n724), .Y(n688) );
  NAND2X1 U724 ( .A(n740), .B(n756), .Y(n748) );
  CLKBUFX3 U725 ( .A(a_11_), .Y(n31) );
  NAND2X1 U726 ( .A(n744), .B(n760), .Y(n752) );
  XNOR2X1 U727 ( .A(n25), .B(n729), .Y(n639) );
  XNOR2X1 U728 ( .A(n728), .B(n25), .Y(n638) );
  CLKINVX1 U729 ( .A(n200), .Y(n198) );
  XNOR2X1 U730 ( .A(n728), .B(n19), .Y(n656) );
  CLKBUFX3 U731 ( .A(a_13_), .Y(n37) );
  CLKBUFX3 U732 ( .A(b_16_), .Y(n721) );
  OAI22X1 U733 ( .A0(n577), .A1(n46), .B0(n48), .B1(n578), .Y(n251) );
  AOI21X1 U734 ( .A0(n113), .A1(n848), .B0(n110), .Y(n108) );
  OAI21X1 U735 ( .A0(n108), .A1(n106), .B0(n107), .Y(n105) );
  OAI21X1 U736 ( .A0(n100), .A1(n98), .B0(n99), .Y(n97) );
  CLKINVX1 U737 ( .A(n120), .Y(n118) );
  AOI21X1 U738 ( .A0(n129), .A1(n844), .B0(n126), .Y(n124) );
  NAND2X1 U739 ( .A(n313), .B(n321), .Y(n131) );
  NOR2X1 U740 ( .A(n313), .B(n321), .Y(n130) );
  OAI21X1 U741 ( .A0(n147), .A1(n145), .B0(n146), .Y(n144) );
  XNOR2X1 U742 ( .A(n735), .B(n43), .Y(n591) );
  OR2X2 U743 ( .A(n393), .B(n400), .Y(n839) );
  INVXL U744 ( .A(a_0_), .Y(n761) );
  OR2X1 U745 ( .A(n419), .B(n423), .Y(n840) );
  NAND2XL U746 ( .A(n754), .B(n738), .Y(n746) );
  BUFX4 U747 ( .A(n746), .Y(n48) );
  OR2X1 U748 ( .A(n322), .B(n332), .Y(n841) );
  XNOR2X2 U749 ( .A(a_11_), .B(a_12_), .Y(n755) );
  OR2X2 U750 ( .A(n401), .B(n406), .Y(n842) );
  OR2X1 U751 ( .A(n424), .B(n425), .Y(n843) );
  OR2X1 U752 ( .A(n312), .B(n303), .Y(n844) );
  OR2X1 U753 ( .A(n432), .B(n574), .Y(n845) );
  OR2X1 U754 ( .A(n426), .B(n429), .Y(n846) );
  OR2X1 U755 ( .A(n294), .B(n287), .Y(n847) );
  OR2X1 U756 ( .A(n274), .B(n280), .Y(n848) );
  OR2X1 U757 ( .A(n268), .B(n264), .Y(n849) );
  OR2X1 U758 ( .A(n256), .B(n260), .Y(n850) );
  OR2X1 U759 ( .A(n253), .B(n252), .Y(n851) );
  BUFX4 U760 ( .A(n750), .Y(n24) );
  BUFX4 U761 ( .A(n749), .Y(n29) );
  BUFX4 U762 ( .A(n753), .Y(n5) );
  XNOR2X1 U763 ( .A(a_13_), .B(a_14_), .Y(n754) );
  CLKBUFX3 U764 ( .A(n747), .Y(n42) );
  CLKBUFX3 U765 ( .A(b_9_), .Y(n728) );
  NOR2BX1 U766 ( .AN(n49), .B(n9), .Y(n559) );
  OAI22X1 U767 ( .A0(n683), .A1(n17), .B0(n682), .B1(n15), .Y(n540) );
  CLKBUFX4 U768 ( .A(a_7_), .Y(n19) );
  OAI22X1 U769 ( .A0(n696), .A1(n11), .B0(n695), .B1(n9), .Y(n553) );
  OAI22X1 U770 ( .A0(n11), .A1(n694), .B0(n693), .B1(n9), .Y(n551) );
  ADDHX2 U771 ( .A(n566), .B(n534), .CO(n397), .S(n398) );
  OAI22X1 U772 ( .A0(n708), .A1(n3), .B0(n753), .B1(n709), .Y(n566) );
  CMPR42X2 U773 ( .A(n553), .B(n420), .C(n537), .D(n416), .ICI(n417), .S(n414), 
        .ICO(n412), .CO(n413) );
  ADDHX1 U774 ( .A(n570), .B(n437), .CO(n420), .S(n421) );
  BUFX4 U775 ( .A(n137), .Y(n852) );
  CLKBUFX4 U776 ( .A(a_5_), .Y(n13) );
  BUFX6 U777 ( .A(n757), .Y(n853) );
  CLKBUFX4 U778 ( .A(a_3_), .Y(n7) );
  CLKBUFX6 U779 ( .A(a_9_), .Y(n25) );
  OAI22X1 U780 ( .A0(n677), .A1(n17), .B0(n676), .B1(n15), .Y(n534) );
  OAI22X1 U781 ( .A0(n681), .A1(n15), .B0(n17), .B1(n682), .Y(n539) );
  CLKINVX1 U782 ( .A(n128), .Y(n126) );
  INVX3 U783 ( .A(n178), .Y(n176) );
  OAI22X1 U784 ( .A0(n702), .A1(n10), .B0(n12), .B1(n768), .Y(n439) );
  OAI22XL U785 ( .A0(n17), .A1(n671), .B0(n670), .B1(n16), .Y(n528) );
  XNOR2XL U786 ( .A(n732), .B(n31), .Y(n624) );
  XNOR2XL U787 ( .A(n7), .B(n725), .Y(n689) );
  XNOR2XL U788 ( .A(n19), .B(n729), .Y(n657) );
  XNOR2X1 U789 ( .A(n129), .B(n62), .Y(product_20_) );
  AOI21X1 U790 ( .A0(n852), .A1(n841), .B0(n134), .Y(n132) );
  CLKBUFX3 U791 ( .A(b_6_), .Y(n731) );
  CLKBUFX2 U792 ( .A(b_7_), .Y(n730) );
  NAND2X1 U793 ( .A(n731), .B(n13), .Y(n855) );
  NAND2X1 U794 ( .A(n854), .B(n767), .Y(n856) );
  NAND2X1 U795 ( .A(n855), .B(n856), .Y(n677) );
  CLKINVX1 U796 ( .A(n731), .Y(n854) );
  OAI22X1 U797 ( .A0(n678), .A1(n17), .B0(n677), .B1(n15), .Y(n535) );
  OR2X8 U798 ( .A(n132), .B(n130), .Y(n857) );
  NAND2X8 U799 ( .A(n857), .B(n131), .Y(n129) );
  OAI21XL U800 ( .A0(n138), .A1(n158), .B0(n139), .Y(n137) );
  NAND2XL U801 ( .A(n140), .B(n148), .Y(n138) );
  CLKBUFX4 U802 ( .A(a_1_), .Y(n1) );
  XNOR2X1 U803 ( .A(n730), .B(n25), .Y(n640) );
  OAI22X1 U804 ( .A0(n648), .A1(n28), .B0(n29), .B1(n765), .Y(n436) );
  XNOR2X1 U805 ( .A(n723), .B(n7), .Y(n687) );
  AOI21X1 U806 ( .A0(n157), .A1(n148), .B0(n149), .Y(n147) );
  INVX1 U807 ( .A(n202), .Y(n201) );
  XNOR2XL U808 ( .A(n730), .B(n13), .Y(n676) );
  XNOR2XL U809 ( .A(n13), .B(n729), .Y(n675) );
  XNOR2XL U810 ( .A(b_9_), .B(n37), .Y(n608) );
  OAI22X1 U811 ( .A0(n701), .A1(n11), .B0(n700), .B1(n9), .Y(n558) );
  OAI22X1 U812 ( .A0(n695), .A1(n11), .B0(n694), .B1(n9), .Y(n552) );
  OAI22X1 U813 ( .A0(n630), .A1(n34), .B0(n36), .B1(n764), .Y(n435) );
  OAI22X1 U814 ( .A0(n629), .A1(n35), .B0(n628), .B1(n33), .Y(n486) );
  CLKBUFX3 U815 ( .A(a_15_), .Y(n43) );
  XNOR2XL U816 ( .A(n733), .B(n31), .Y(n625) );
  OAI21XL U817 ( .A0(n142), .A1(n146), .B0(n143), .Y(n141) );
  CLKBUFX4 U818 ( .A(b_0_), .Y(n49) );
  OAI21X1 U819 ( .A0(n208), .A1(n210), .B0(n209), .Y(n207) );
  NAND2BXL U820 ( .AN(n218), .B(n219), .Y(n81) );
  INVX1 U821 ( .A(n81), .Y(product_1_) );
  CMPR42X1 U822 ( .A(n518), .B(n550), .C(n403), .D(n399), .ICI(n396), .S(n393), 
        .ICO(n391), .CO(n392) );
  NOR2BXL U823 ( .AN(n49), .B(n3), .Y(product_0_) );
  AO21XL U824 ( .A0(n42), .A1(n40), .B0(n595), .Y(n456) );
  XNOR2X1 U825 ( .A(n730), .B(n1), .Y(n712) );
  XNOR2X1 U826 ( .A(n731), .B(n1), .Y(n713) );
  XNOR2X1 U827 ( .A(n7), .B(n722), .Y(n686) );
  XNOR2X1 U828 ( .A(a_7_), .B(a_8_), .Y(n757) );
  INVX3 U829 ( .A(n158), .Y(n157) );
  OAI21X2 U830 ( .A0(n180), .A1(n168), .B0(n169), .Y(n167) );
  NAND2XL U831 ( .A(n238), .B(n162), .Y(n69) );
  AOI21XL U832 ( .A0(n140), .A1(n149), .B0(n141), .Y(n139) );
  CLKBUFX2 U833 ( .A(b_12_), .Y(n725) );
  INVXL U834 ( .A(n180), .Y(n179) );
  NAND2XL U835 ( .A(n234), .B(n143), .Y(n65) );
  NAND2XL U836 ( .A(n236), .B(n151), .Y(n67) );
  NAND2XL U837 ( .A(n839), .B(n173), .Y(n71) );
  XNOR2X1 U838 ( .A(n858), .B(n51), .Y(product_31_) );
  AO21XL U839 ( .A0(n89), .A1(n851), .B0(n86), .Y(n858) );
  INVXL U840 ( .A(n156), .Y(n154) );
  INVXL U841 ( .A(n161), .Y(n238) );
  NOR2X1 U842 ( .A(n355), .B(n365), .Y(n150) );
  NOR2X1 U843 ( .A(n366), .B(n374), .Y(n155) );
  NOR2X1 U844 ( .A(n385), .B(n392), .Y(n164) );
  CLKBUFX2 U845 ( .A(b_14_), .Y(n723) );
  NOR2X1 U846 ( .A(n333), .B(n343), .Y(n142) );
  NOR2X1 U847 ( .A(n344), .B(n354), .Y(n145) );
  NOR2X1 U848 ( .A(n302), .B(n295), .Y(n122) );
  NOR2X1 U849 ( .A(n281), .B(n286), .Y(n114) );
  NOR2X1 U850 ( .A(n269), .B(n273), .Y(n106) );
  NOR2X1 U851 ( .A(n254), .B(n255), .Y(n90) );
  CLKBUFX2 U852 ( .A(b_8_), .Y(n729) );
  NOR2BXL U853 ( .AN(n49), .B(n33), .Y(n487) );
  NOR2X1 U854 ( .A(n414), .B(n418), .Y(n186) );
  NOR2X1 U855 ( .A(n575), .B(n559), .Y(n216) );
  NOR2XL U856 ( .A(n838), .B(n440), .Y(n218) );
  NOR2X1 U857 ( .A(n430), .B(n431), .Y(n208) );
  CMPR32X2 U858 ( .A(n572), .B(n556), .C(n428), .CO(n425), .S(n426) );
  XNOR2XL U859 ( .A(b_9_), .B(n43), .Y(n590) );
  XNOR2XL U860 ( .A(n49), .B(n43), .Y(n593) );
  NAND2BXL U861 ( .AN(n49), .B(n43), .Y(n594) );
  XNOR2XL U862 ( .A(n733), .B(n43), .Y(n589) );
  XNOR2XL U863 ( .A(n732), .B(n43), .Y(n588) );
  XNOR2XL U864 ( .A(n731), .B(n43), .Y(n587) );
  XNOR2XL U865 ( .A(n730), .B(n43), .Y(n586) );
  XNOR2XL U866 ( .A(n728), .B(n43), .Y(n584) );
  XNOR2XL U867 ( .A(n729), .B(n43), .Y(n585) );
  OAI22XL U868 ( .A0(n35), .A1(n622), .B0(n621), .B1(n33), .Y(n329) );
  AO21XL U869 ( .A0(n749), .A1(n28), .B0(n631), .Y(n488) );
  XNOR2XL U870 ( .A(n726), .B(n43), .Y(n582) );
  XNOR2XL U871 ( .A(n725), .B(n43), .Y(n581) );
  XNOR2XL U872 ( .A(n43), .B(n722), .Y(n583) );
  NOR2X1 U873 ( .A(n261), .B(n263), .Y(n98) );
  ADDFXL U874 ( .A(n258), .B(n259), .CI(n457), .CO(n255), .S(n256) );
  XNOR2XL U875 ( .A(n723), .B(n43), .Y(n579) );
  ADDFXL U876 ( .A(n442), .B(n257), .CI(n456), .CO(n253), .S(n254) );
  AO21XL U877 ( .A0(n48), .A1(n46), .B0(n577), .Y(n441) );
  XNOR2XL U878 ( .A(n49), .B(n7), .Y(n701) );
  XNOR2XL U879 ( .A(n735), .B(n13), .Y(n681) );
  XNOR2XL U880 ( .A(n732), .B(n7), .Y(n696) );
  XNOR2XL U881 ( .A(n733), .B(n1), .Y(n715) );
  XNOR2XL U882 ( .A(n733), .B(n7), .Y(n697) );
  XNOR2XL U883 ( .A(n732), .B(n1), .Y(n714) );
  XNOR2XL U884 ( .A(n735), .B(n25), .Y(n645) );
  XNOR2XL U885 ( .A(n731), .B(n19), .Y(n659) );
  XNOR2XL U886 ( .A(n735), .B(n31), .Y(n627) );
  XNOR2XL U887 ( .A(n732), .B(n19), .Y(n660) );
  XNOR2XL U888 ( .A(n732), .B(n25), .Y(n642) );
  XNOR2XL U889 ( .A(n733), .B(n19), .Y(n661) );
  XNOR2XL U890 ( .A(n733), .B(n25), .Y(n643) );
  XNOR2XL U891 ( .A(b_9_), .B(n13), .Y(n680) );
  XNOR2XL U892 ( .A(b_3_), .B(n7), .Y(n698) );
  XNOR2XL U893 ( .A(n728), .B(n7), .Y(n692) );
  XNOR2XL U894 ( .A(b_9_), .B(n31), .Y(n626) );
  XNOR2XL U895 ( .A(n7), .B(n729), .Y(n693) );
  CLKBUFX2 U896 ( .A(n758), .Y(n22) );
  ADDFX2 U897 ( .A(n382), .B(n516), .CI(n434), .CO(n379), .S(n380) );
  OAI22X1 U898 ( .A0(n612), .A1(n40), .B0(n42), .B1(n763), .Y(n434) );
  CLKBUFX2 U899 ( .A(n758), .Y(n21) );
  XNOR2XL U900 ( .A(n49), .B(n13), .Y(n683) );
  XNOR2XL U901 ( .A(n49), .B(n19), .Y(n665) );
  XNOR2XL U902 ( .A(n49), .B(n31), .Y(n629) );
  XNOR2XL U903 ( .A(n49), .B(n37), .Y(n611) );
  NAND2BXL U904 ( .AN(n49), .B(n1), .Y(n720) );
  NAND2BXL U905 ( .AN(n49), .B(n25), .Y(n648) );
  NAND2BXL U906 ( .AN(n49), .B(n19), .Y(n666) );
  NAND2BXL U907 ( .AN(n49), .B(n7), .Y(n702) );
  NAND2BXL U908 ( .AN(n49), .B(n13), .Y(n684) );
  NAND2BXL U909 ( .AN(n49), .B(n31), .Y(n630) );
  NAND2BXL U910 ( .AN(n49), .B(n37), .Y(n612) );
  CMPR32X2 U911 ( .A(n541), .B(n557), .C(n573), .CO(n429), .S(n430) );
  NOR2BXL U912 ( .AN(n49), .B(n15), .Y(n541) );
  XNOR2XL U913 ( .A(n13), .B(n725), .Y(n671) );
  XNOR2XL U914 ( .A(n730), .B(n19), .Y(n658) );
  XNOR2XL U915 ( .A(n735), .B(n37), .Y(n609) );
  XNOR2XL U916 ( .A(n731), .B(n25), .Y(n641) );
  XNOR2XL U917 ( .A(n731), .B(n31), .Y(n623) );
  XNOR2XL U918 ( .A(n733), .B(n37), .Y(n607) );
  XNOR2XL U919 ( .A(n732), .B(n37), .Y(n606) );
  XNOR2XL U920 ( .A(n728), .B(n13), .Y(n674) );
  XNOR2XL U921 ( .A(n726), .B(n13), .Y(n672) );
  XNOR2XL U922 ( .A(n726), .B(n19), .Y(n654) );
  XNOR2XL U923 ( .A(n19), .B(n725), .Y(n653) );
  XNOR2XL U924 ( .A(n721), .B(n7), .Y(n685) );
  XNOR2XL U925 ( .A(n13), .B(b_10_), .Y(n673) );
  XNOR2XL U926 ( .A(n19), .B(n722), .Y(n655) );
  XNOR2XL U927 ( .A(n723), .B(n31), .Y(n615) );
  XNOR2XL U928 ( .A(n31), .B(n729), .Y(n621) );
  XNOR2XL U929 ( .A(n723), .B(n13), .Y(n669) );
  XNOR2XL U930 ( .A(n730), .B(n37), .Y(n604) );
  XNOR2XL U931 ( .A(n723), .B(n19), .Y(n651) );
  XNOR2XL U932 ( .A(n723), .B(n25), .Y(n633) );
  XNOR2XL U933 ( .A(n731), .B(n37), .Y(n605) );
  XNOR2XL U934 ( .A(n728), .B(n31), .Y(n620) );
  XNOR2XL U935 ( .A(n726), .B(n25), .Y(n636) );
  XNOR2XL U936 ( .A(n726), .B(n37), .Y(n600) );
  XNOR2XL U937 ( .A(n728), .B(n37), .Y(n602) );
  XNOR2XL U938 ( .A(n726), .B(n31), .Y(n618) );
  XNOR2XL U939 ( .A(n25), .B(n725), .Y(n635) );
  XNOR2XL U940 ( .A(n37), .B(n725), .Y(n599) );
  XNOR2XL U941 ( .A(n31), .B(n725), .Y(n617) );
  XNOR2XL U942 ( .A(n721), .B(n13), .Y(n667) );
  XNOR2XL U943 ( .A(n721), .B(n25), .Y(n631) );
  XNOR2XL U944 ( .A(n721), .B(n19), .Y(n649) );
  XNOR2XL U945 ( .A(n37), .B(n729), .Y(n603) );
  XNOR2XL U946 ( .A(n13), .B(n722), .Y(n668) );
  XNOR2XL U947 ( .A(n25), .B(n722), .Y(n637) );
  XNOR2XL U948 ( .A(n19), .B(n722), .Y(n650) );
  XNOR2XL U949 ( .A(n25), .B(n722), .Y(n632) );
  XNOR2XL U950 ( .A(n37), .B(n722), .Y(n601) );
  XNOR2XL U951 ( .A(n31), .B(n722), .Y(n619) );
  OAI22XL U952 ( .A0(n36), .A1(n616), .B0(n615), .B1(n34), .Y(n277) );
  XNOR2XL U953 ( .A(n723), .B(n37), .Y(n597) );
  XNOR2XL U954 ( .A(n721), .B(n37), .Y(n595) );
  XNOR2XL U955 ( .A(n721), .B(n31), .Y(n613) );
  XNOR2XL U956 ( .A(n31), .B(n722), .Y(n614) );
  OAI22XL U957 ( .A0(n42), .A1(n598), .B0(n597), .B1(n40), .Y(n265) );
  AO21XL U958 ( .A0(n36), .A1(n34), .B0(n613), .Y(n472) );
  XNOR2XL U959 ( .A(n37), .B(n722), .Y(n596) );
  OAI22XL U960 ( .A0(n579), .A1(n46), .B0(n48), .B1(n580), .Y(n257) );
  XNOR2X1 U961 ( .A(a_3_), .B(a_4_), .Y(n759) );
  XNOR2X1 U962 ( .A(a_1_), .B(a_2_), .Y(n760) );
  XNOR2X1 U963 ( .A(a_9_), .B(a_10_), .Y(n756) );
  XNOR2XL U964 ( .A(n13), .B(n724), .Y(n670) );
  XNOR2XL U965 ( .A(n19), .B(n724), .Y(n652) );
  XNOR2XL U966 ( .A(n25), .B(n724), .Y(n634) );
  XNOR2XL U967 ( .A(n43), .B(n724), .Y(n580) );
  CLKBUFX2 U968 ( .A(b_13_), .Y(n724) );
  CLKBUFX3 U969 ( .A(b_11_), .Y(n726) );
  XNOR2X1 U970 ( .A(n179), .B(n72), .Y(product_10_) );
  NAND2X1 U971 ( .A(n842), .B(n178), .Y(n72) );
  NAND2X1 U972 ( .A(n839), .B(n842), .Y(n168) );
  AOI21X1 U973 ( .A0(n839), .A1(n176), .B0(n171), .Y(n169) );
  AOI21X1 U974 ( .A0(n167), .A1(n159), .B0(n160), .Y(n158) );
  OAI21XL U975 ( .A0(n161), .A1(n165), .B0(n162), .Y(n160) );
  NOR2X1 U976 ( .A(n164), .B(n161), .Y(n159) );
  CLKINVX1 U977 ( .A(n136), .Y(n134) );
  CLKINVX1 U978 ( .A(n112), .Y(n110) );
  AOI21X1 U979 ( .A0(n105), .A1(n849), .B0(n102), .Y(n100) );
  CLKINVX1 U980 ( .A(n104), .Y(n102) );
  OAI21X1 U981 ( .A0(n150), .A1(n156), .B0(n151), .Y(n149) );
  OAI21X1 U982 ( .A0(n124), .A1(n122), .B0(n123), .Y(n121) );
  CLKBUFX3 U983 ( .A(b_4_), .Y(n733) );
  CLKBUFX3 U984 ( .A(b_5_), .Y(n732) );
  NOR2X1 U985 ( .A(n142), .B(n145), .Y(n140) );
  NOR2X1 U986 ( .A(n155), .B(n150), .Y(n148) );
  CLKINVX1 U987 ( .A(n189), .Y(n188) );
  XNOR2X1 U988 ( .A(n157), .B(n68), .Y(product_14_) );
  NAND2X1 U989 ( .A(n153), .B(n156), .Y(n68) );
  XNOR2X1 U990 ( .A(n144), .B(n65), .Y(product_17_) );
  XNOR2X1 U991 ( .A(n163), .B(n69), .Y(product_13_) );
  XNOR2X1 U992 ( .A(n89), .B(n52), .Y(product_30_) );
  NAND2X1 U993 ( .A(n851), .B(n88), .Y(n52) );
  XNOR2X1 U994 ( .A(n105), .B(n56), .Y(product_26_) );
  NAND2X1 U995 ( .A(n849), .B(n104), .Y(n56) );
  XNOR2X1 U996 ( .A(n113), .B(n58), .Y(product_24_) );
  NAND2X1 U997 ( .A(n848), .B(n112), .Y(n58) );
  XNOR2X1 U998 ( .A(n121), .B(n60), .Y(product_22_) );
  NAND2X1 U999 ( .A(n847), .B(n120), .Y(n60) );
  NAND2X1 U1000 ( .A(n844), .B(n128), .Y(n62) );
  XNOR2X1 U1001 ( .A(n852), .B(n64), .Y(product_18_) );
  NAND2X1 U1002 ( .A(n841), .B(n136), .Y(n64) );
  CLKINVX1 U1003 ( .A(n155), .Y(n153) );
  CLKINVX1 U1004 ( .A(n173), .Y(n171) );
  XOR2X1 U1005 ( .A(n174), .B(n71), .Y(product_11_) );
  AOI21X1 U1006 ( .A0(n179), .A1(n842), .B0(n176), .Y(n174) );
  XOR2X1 U1007 ( .A(n166), .B(n70), .Y(product_12_) );
  NAND2X1 U1008 ( .A(n239), .B(n165), .Y(n70) );
  CLKINVX1 U1009 ( .A(n164), .Y(n239) );
  XOR2X1 U1010 ( .A(n152), .B(n67), .Y(product_15_) );
  AOI21X1 U1011 ( .A0(n157), .A1(n153), .B0(n154), .Y(n152) );
  NAND2X1 U1012 ( .A(n859), .B(n83), .Y(n51) );
  XOR2X1 U1013 ( .A(n147), .B(n66), .Y(product_16_) );
  NAND2X1 U1014 ( .A(n235), .B(n146), .Y(n66) );
  CLKINVX1 U1015 ( .A(n145), .Y(n235) );
  XOR2X1 U1016 ( .A(n92), .B(n53), .Y(product_29_) );
  NAND2X1 U1017 ( .A(n222), .B(n91), .Y(n53) );
  CLKINVX1 U1018 ( .A(n90), .Y(n222) );
  XOR2X1 U1019 ( .A(n108), .B(n57), .Y(product_25_) );
  NAND2X1 U1020 ( .A(n226), .B(n107), .Y(n57) );
  CLKINVX1 U1021 ( .A(n106), .Y(n226) );
  XOR2X1 U1022 ( .A(n116), .B(n59), .Y(product_23_) );
  NAND2X1 U1023 ( .A(n228), .B(n115), .Y(n59) );
  CLKINVX1 U1024 ( .A(n114), .Y(n228) );
  XOR2X1 U1025 ( .A(n124), .B(n61), .Y(product_21_) );
  NAND2X1 U1026 ( .A(n230), .B(n123), .Y(n61) );
  CLKINVX1 U1027 ( .A(n122), .Y(n230) );
  XOR2X1 U1028 ( .A(n132), .B(n63), .Y(product_19_) );
  NAND2X1 U1029 ( .A(n232), .B(n131), .Y(n63) );
  CLKINVX1 U1030 ( .A(n130), .Y(n232) );
  CLKINVX1 U1031 ( .A(n183), .Y(n242) );
  CLKINVX1 U1032 ( .A(n142), .Y(n234) );
  CLKINVX1 U1033 ( .A(n150), .Y(n236) );
  CLKINVX1 U1034 ( .A(n88), .Y(n86) );
  CMPR42X1 U1035 ( .A(n334), .B(n338), .C(n335), .D(n325), .ICI(n331), .S(n322), .ICO(n320), .CO(n321) );
  XNOR2X1 U1036 ( .A(n79), .B(n215), .Y(product_3_) );
  NAND2X1 U1037 ( .A(n845), .B(n214), .Y(n79) );
  AOI21X1 U1038 ( .A0(n181), .A1(n189), .B0(n182), .Y(n180) );
  NOR2X1 U1039 ( .A(n183), .B(n186), .Y(n181) );
  OAI21XL U1040 ( .A0(n183), .A1(n187), .B0(n184), .Y(n182) );
  NAND2X1 U1041 ( .A(n840), .B(n843), .Y(n190) );
  AOI21X1 U1042 ( .A0(n840), .A1(n198), .B0(n193), .Y(n191) );
  AOI21X1 U1043 ( .A0(n207), .A1(n846), .B0(n204), .Y(n202) );
  CLKINVX1 U1044 ( .A(n206), .Y(n204) );
  NOR2X2 U1045 ( .A(n375), .B(n384), .Y(n161) );
  CLKINVX1 U1046 ( .A(n96), .Y(n94) );
  AOI21X1 U1047 ( .A0(n215), .A1(n845), .B0(n212), .Y(n210) );
  CLKINVX1 U1048 ( .A(n214), .Y(n212) );
  OAI21X1 U1049 ( .A0(n216), .A1(n219), .B0(n217), .Y(n215) );
  NAND2X1 U1050 ( .A(n366), .B(n374), .Y(n156) );
  NAND2X1 U1051 ( .A(n385), .B(n392), .Y(n165) );
  NAND2X1 U1052 ( .A(n344), .B(n354), .Y(n146) );
  NAND2X1 U1053 ( .A(n312), .B(n303), .Y(n128) );
  NAND2X1 U1054 ( .A(n393), .B(n400), .Y(n173) );
  NAND2X1 U1055 ( .A(n401), .B(n406), .Y(n178) );
  NAND2X1 U1056 ( .A(n322), .B(n332), .Y(n136) );
  NAND2X1 U1057 ( .A(n407), .B(n413), .Y(n184) );
  NAND2X1 U1058 ( .A(n375), .B(n384), .Y(n162) );
  NAND2X1 U1059 ( .A(n355), .B(n365), .Y(n151) );
  NAND2X1 U1060 ( .A(n333), .B(n343), .Y(n143) );
  XOR2X1 U1061 ( .A(n78), .B(n210), .Y(product_4_) );
  NAND2X1 U1062 ( .A(n247), .B(n209), .Y(n78) );
  CLKINVX1 U1063 ( .A(n208), .Y(n247) );
  XOR2X1 U1064 ( .A(n80), .B(n219), .Y(product_2_) );
  NAND2X1 U1065 ( .A(n249), .B(n217), .Y(n80) );
  CLKINVX1 U1066 ( .A(n216), .Y(n249) );
  XNOR2X1 U1067 ( .A(n201), .B(n76), .Y(product_6_) );
  NAND2X1 U1068 ( .A(n843), .B(n200), .Y(n76) );
  CLKINVX1 U1069 ( .A(n329), .Y(n330) );
  NAND2X1 U1070 ( .A(n242), .B(n184), .Y(n73) );
  XNOR2X1 U1071 ( .A(n97), .B(n54), .Y(product_28_) );
  NAND2X1 U1072 ( .A(n850), .B(n96), .Y(n54) );
  XNOR2X1 U1073 ( .A(n207), .B(n77), .Y(product_5_) );
  NAND2X1 U1074 ( .A(n846), .B(n206), .Y(n77) );
  CLKINVX1 U1075 ( .A(n195), .Y(n193) );
  XOR2X1 U1076 ( .A(n188), .B(n74), .Y(product_8_) );
  NAND2X1 U1077 ( .A(n243), .B(n187), .Y(n74) );
  CLKINVX1 U1078 ( .A(n186), .Y(n243) );
  XOR2X1 U1079 ( .A(n196), .B(n75), .Y(product_7_) );
  NAND2X1 U1080 ( .A(n840), .B(n195), .Y(n75) );
  AOI21X1 U1081 ( .A0(n201), .A1(n843), .B0(n198), .Y(n196) );
  XOR2X1 U1082 ( .A(n100), .B(n55), .Y(product_27_) );
  NAND2X1 U1083 ( .A(n224), .B(n99), .Y(n55) );
  CLKINVX1 U1084 ( .A(n98), .Y(n224) );
  NAND2X1 U1085 ( .A(n294), .B(n287), .Y(n120) );
  NAND2X1 U1086 ( .A(n268), .B(n264), .Y(n104) );
  NAND2X1 U1087 ( .A(n274), .B(n280), .Y(n112) );
  NAND2X1 U1088 ( .A(n302), .B(n295), .Y(n123) );
  NAND2X1 U1089 ( .A(n281), .B(n286), .Y(n115) );
  NAND2X1 U1090 ( .A(n269), .B(n273), .Y(n107) );
  NAND2X1 U1091 ( .A(n441), .B(n251), .Y(n83) );
  NAND2X1 U1092 ( .A(n253), .B(n252), .Y(n88) );
  CLKINVX1 U1093 ( .A(n251), .Y(n252) );
  NAND2X1 U1094 ( .A(n254), .B(n255), .Y(n91) );
  OR2X1 U1095 ( .A(n441), .B(n251), .Y(n859) );
  OAI22XL U1096 ( .A0(n747), .A1(n604), .B0(n603), .B1(n755), .Y(n309) );
  OAI22XL U1097 ( .A0(n661), .A1(n24), .B0(n660), .B1(n21), .Y(n518) );
  OAI22XL U1098 ( .A0(n692), .A1(n10), .B0(n11), .B1(n693), .Y(n550) );
  OAI22XL U1099 ( .A0(n710), .A1(n3), .B0(n5), .B1(n711), .Y(n568) );
  OAI22XL U1100 ( .A0(n656), .A1(n21), .B0(n663), .B1(n24), .Y(n520) );
  OAI22XL U1101 ( .A0(n680), .A1(n17), .B0(n679), .B1(n15), .Y(n537) );
  CMPR42X1 U1102 ( .A(n532), .B(n380), .C(n387), .D(n378), .ICI(n383), .S(n375), .ICO(n373), .CO(n374) );
  OAI22XL U1103 ( .A0(n674), .A1(n16), .B0(n17), .B1(n675), .Y(n532) );
  CMPR42X1 U1104 ( .A(n390), .B(n549), .C(n395), .D(n391), .ICI(n388), .S(n385), .ICO(n383), .CO(n384) );
  OAI22XL U1105 ( .A0(n692), .A1(n12), .B0(n691), .B1(n10), .Y(n549) );
  CMPR42X1 U1106 ( .A(n371), .B(n361), .C(n368), .D(n358), .ICI(n364), .S(n355), .ICO(n353), .CO(n354) );
  CMPR42X1 U1107 ( .A(n379), .B(n372), .C(n377), .D(n369), .ICI(n373), .S(n366), .ICO(n364), .CO(n365) );
  CMPR42X1 U1108 ( .A(n339), .B(n560), .C(n346), .D(n342), .ICI(n336), .S(n333), .ICO(n331), .CO(n332) );
  AO21X1 U1109 ( .A0(n753), .A1(n3), .B0(n703), .Y(n560) );
  CMPR42X1 U1110 ( .A(n350), .B(n561), .C(n357), .D(n353), .ICI(n347), .S(n344), .ICO(n342), .CO(n343) );
  OAI22XL U1111 ( .A0(n703), .A1(n3), .B0(n753), .B1(n704), .Y(n561) );
  CMPR42X1 U1112 ( .A(n323), .B(n542), .C(n324), .D(n316), .ICI(n320), .S(n313), .ICO(n311), .CO(n312) );
  AO21X1 U1113 ( .A0(n12), .A1(n10), .B0(n685), .Y(n542) );
  CMPR42X1 U1114 ( .A(n314), .B(n525), .C(n306), .D(n315), .ICI(n311), .S(n303), .ICO(n301), .CO(n302) );
  OAI22XL U1115 ( .A0(n667), .A1(n16), .B0(n17), .B1(n668), .Y(n525) );
  OAI22XL U1116 ( .A0(n12), .A1(n687), .B0(n686), .B1(n10), .Y(n544) );
  XNOR2X1 U1117 ( .A(n544), .B(n528), .Y(n341) );
  OAI22XL U1118 ( .A0(n608), .A1(n40), .B0(n609), .B1(n747), .Y(n468) );
  OAI22XL U1119 ( .A0(n626), .A1(n35), .B0(n625), .B1(n33), .Y(n483) );
  OAI22XL U1120 ( .A0(n690), .A1(n12), .B0(n689), .B1(n10), .Y(n547) );
  OAI22XL U1121 ( .A0(n698), .A1(n11), .B0(n697), .B1(n9), .Y(n555) );
  OAI22XL U1122 ( .A0(n715), .A1(n5), .B0(n714), .B1(n3), .Y(n572) );
  OAI22XL U1123 ( .A0(n698), .A1(n9), .B0(n699), .B1(n11), .Y(n556) );
  NAND2X1 U1124 ( .A(n414), .B(n418), .Y(n187) );
  CMPR42X1 U1125 ( .A(n512), .B(n351), .C(n341), .D(n480), .ICI(n466), .S(n339), .ICO(n337), .CO(n338) );
  OAI22XL U1126 ( .A0(n607), .A1(n747), .B0(n606), .B1(n40), .Y(n466) );
  OAI22XL U1127 ( .A0(n654), .A1(n22), .B0(n24), .B1(n655), .Y(n512) );
  OAI22XL U1128 ( .A0(n623), .A1(n35), .B0(n622), .B1(n33), .Y(n480) );
  NAND2X1 U1129 ( .A(n419), .B(n423), .Y(n195) );
  CMPR42X1 U1130 ( .A(n317), .B(n308), .C(n449), .D(n478), .ICI(n318), .S(n306), .ICO(n304), .CO(n305) );
  OAI22XL U1131 ( .A0(n588), .A1(n48), .B0(n587), .B1(n46), .Y(n449) );
  OAI22XL U1132 ( .A0(n620), .A1(n36), .B0(n619), .B1(n34), .Y(n478) );
  NAND2X1 U1133 ( .A(n424), .B(n425), .Y(n200) );
  NAND2X1 U1134 ( .A(n575), .B(n559), .Y(n217) );
  NAND2X1 U1135 ( .A(n432), .B(n574), .Y(n214) );
  CMPR42X1 U1136 ( .A(n481), .B(n513), .C(n467), .D(n356), .ICI(n360), .S(n347), .ICO(n345), .CO(n346) );
  OAI22XL U1137 ( .A0(n624), .A1(n35), .B0(n623), .B1(n33), .Y(n481) );
  OAI22XL U1138 ( .A0(n608), .A1(n747), .B0(n607), .B1(n40), .Y(n467) );
  OAI22XL U1139 ( .A0(n656), .A1(n24), .B0(n655), .B1(n22), .Y(n513) );
  NAND2X1 U1140 ( .A(n426), .B(n429), .Y(n206) );
  CMPR42X1 U1141 ( .A(n433), .B(n482), .C(n468), .D(n514), .ICI(n367), .S(n358), .ICO(n356), .CO(n357) );
  OAI22XL U1142 ( .A0(n625), .A1(n35), .B0(n624), .B1(n33), .Y(n482) );
  OAI22XL U1143 ( .A0(n594), .A1(n46), .B0(n48), .B1(n762), .Y(n433) );
  OAI22XL U1144 ( .A0(n656), .A1(n22), .B0(n750), .B1(n657), .Y(n514) );
  CMPR42X1 U1145 ( .A(n527), .B(n511), .C(n330), .D(n340), .ICI(n465), .S(n328), .ICO(n326), .CO(n327) );
  OAI22XL U1146 ( .A0(n606), .A1(n42), .B0(n605), .B1(n755), .Y(n465) );
  OAI22XL U1147 ( .A0(n654), .A1(n24), .B0(n653), .B1(n22), .Y(n511) );
  OR2X1 U1148 ( .A(n544), .B(n528), .Y(n340) );
  CMPR42X1 U1149 ( .A(n326), .B(n464), .C(n479), .D(n327), .ICI(n319), .S(n316), .ICO(n314), .CO(n315) );
  OAI22XL U1150 ( .A0(n605), .A1(n42), .B0(n604), .B1(n755), .Y(n464) );
  OAI22XL U1151 ( .A0(n620), .A1(n34), .B0(n35), .B1(n621), .Y(n479) );
  CMPR42X1 U1152 ( .A(n337), .B(n451), .C(n495), .D(n328), .ICI(n543), .S(n325), .ICO(n323), .CO(n324) );
  OAI22XL U1153 ( .A0(n685), .A1(n10), .B0(n12), .B1(n686), .Y(n543) );
  OAI22XL U1154 ( .A0(n638), .A1(n29), .B0(n637), .B1(n28), .Y(n495) );
  OAI22XL U1155 ( .A0(n590), .A1(n48), .B0(n589), .B1(n46), .Y(n451) );
  CMPR42X1 U1156 ( .A(n567), .B(n519), .C(n408), .D(n405), .ICI(n404), .S(n401), .ICO(n399), .CO(n400) );
  OAI22XL U1157 ( .A0(n656), .A1(n24), .B0(n661), .B1(n21), .Y(n519) );
  OAI22XL U1158 ( .A0(n710), .A1(n753), .B0(n709), .B1(n3), .Y(n567) );
  NAND2X1 U1159 ( .A(n430), .B(n431), .Y(n209) );
  CMPR42X1 U1160 ( .A(n348), .B(n496), .C(n452), .D(n349), .ICI(n345), .S(n336), .ICO(n334), .CO(n335) );
  OAI22XL U1161 ( .A0(n590), .A1(n46), .B0(n591), .B1(n48), .Y(n452) );
  OAI22XL U1162 ( .A0(n638), .A1(n28), .B0(n29), .B1(n639), .Y(n496) );
  CMPR42X1 U1163 ( .A(n510), .B(n329), .C(n526), .D(n494), .ICI(n450), .S(n319), .ICO(n317), .CO(n318) );
  OAI22XL U1164 ( .A0(n636), .A1(n28), .B0(n29), .B1(n637), .Y(n494) );
  OAI22XL U1165 ( .A0(n17), .A1(n669), .B0(n668), .B1(n16), .Y(n526) );
  OAI22XL U1166 ( .A0(n589), .A1(n48), .B0(n588), .B1(n46), .Y(n450) );
  ADDFXL U1167 ( .A(n533), .B(n565), .CI(n471), .CO(n389), .S(n390) );
  OAI22XL U1168 ( .A0(n708), .A1(n5), .B0(n707), .B1(n3), .Y(n565) );
  NOR2BX1 U1169 ( .AN(n49), .B(n40), .Y(n471) );
  OAI22XL U1170 ( .A0(n586), .A1(n48), .B0(n46), .B1(n585), .Y(n291) );
  CMPR42X1 U1171 ( .A(n276), .B(n446), .C(n283), .D(n489), .ICI(n279), .S(n274), .ICO(n272), .CO(n273) );
  OAI22XL U1172 ( .A0(n584), .A1(n48), .B0(n46), .B1(n583), .Y(n446) );
  OAI22XL U1173 ( .A0(n631), .A1(n28), .B0(n29), .B1(n632), .Y(n489) );
  CMPR42X1 U1174 ( .A(n445), .B(n271), .C(n275), .D(n272), .ICI(n488), .S(n269), .ICO(n267), .CO(n268) );
  OAI22XL U1175 ( .A0(n582), .A1(n46), .B0(n48), .B1(n583), .Y(n445) );
  CMPR42X1 U1176 ( .A(n447), .B(n284), .C(n289), .D(n506), .ICI(n285), .S(n281), .ICO(n279), .CO(n280) );
  OAI22XL U1177 ( .A0(n584), .A1(n46), .B0(n48), .B1(n585), .Y(n447) );
  AO21X1 U1178 ( .A0(n24), .A1(n22), .B0(n649), .Y(n506) );
  CMPR42X1 U1179 ( .A(n444), .B(n266), .C(n270), .D(n267), .ICI(n473), .S(n264), .ICO(n262), .CO(n263) );
  OAI22XL U1180 ( .A0(n582), .A1(n48), .B0(n46), .B1(n581), .Y(n444) );
  CLKINVX1 U1181 ( .A(n265), .Y(n266) );
  OAI22XL U1182 ( .A0(n613), .A1(n34), .B0(n36), .B1(n614), .Y(n473) );
  CMPR42X1 U1183 ( .A(n462), .B(n290), .C(n507), .D(n297), .ICI(n293), .S(n287), .ICO(n285), .CO(n286) );
  OAI22XL U1184 ( .A0(n602), .A1(n42), .B0(n601), .B1(n40), .Y(n462) );
  OAI22XL U1185 ( .A0(n649), .A1(n22), .B0(n24), .B1(n650), .Y(n507) );
  CMPR42X1 U1186 ( .A(n304), .B(n524), .C(n298), .D(n305), .ICI(n301), .S(n295), .ICO(n293), .CO(n294) );
  AO21X1 U1187 ( .A0(n17), .A1(n16), .B0(n667), .Y(n524) );
  CLKBUFX3 U1188 ( .A(b_15_), .Y(n722) );
  CMPR42X1 U1189 ( .A(n477), .B(n300), .C(n307), .D(n448), .ICI(n463), .S(n298), .ICO(n296), .CO(n297) );
  OAI22XL U1190 ( .A0(n618), .A1(n34), .B0(n36), .B1(n619), .Y(n477) );
  OAI22XL U1191 ( .A0(n602), .A1(n40), .B0(n42), .B1(n603), .Y(n463) );
  OAI22XL U1192 ( .A0(n587), .A1(n48), .B0(n586), .B1(n46), .Y(n448) );
  ADDFXL U1193 ( .A(n460), .B(n278), .CI(n282), .CO(n275), .S(n276) );
  OAI22XL U1194 ( .A0(n600), .A1(n42), .B0(n599), .B1(n40), .Y(n460) );
  CLKINVX1 U1195 ( .A(n277), .Y(n278) );
  CLKINVX1 U1196 ( .A(n43), .Y(n762) );
  XNOR2X1 U1197 ( .A(n721), .B(n43), .Y(n577) );
  CLKINVX1 U1198 ( .A(n257), .Y(n258) );
  OAI22XL U1199 ( .A0(n595), .A1(n40), .B0(n42), .B1(n596), .Y(n457) );
  OAI22XL U1200 ( .A0(n579), .A1(n48), .B0(n46), .B1(n578), .Y(n442) );
  NAND2X1 U1201 ( .A(n256), .B(n260), .Y(n96) );
  NAND2X1 U1202 ( .A(n261), .B(n263), .Y(n99) );
  XNOR2X1 U1203 ( .A(n43), .B(n722), .Y(n578) );
  XNOR2X1 U1204 ( .A(n49), .B(n1), .Y(n719) );
  OAI22X1 U1205 ( .A0(n717), .A1(n3), .B0(n5), .B1(n718), .Y(n575) );
  CLKINVX1 U1206 ( .A(n1), .Y(n769) );
  OAI22XL U1207 ( .A0(n665), .A1(n24), .B0(n664), .B1(n21), .Y(n522) );
  OAI22XL U1208 ( .A0(n680), .A1(n15), .B0(n681), .B1(n17), .Y(n538) );
  CMPR42X1 U1209 ( .A(n523), .B(n539), .C(n571), .D(n555), .ICI(n427), .S(n424), .ICO(n422), .CO(n423) );
  OAI22XL U1210 ( .A0(n714), .A1(n5), .B0(n713), .B1(n3), .Y(n571) );
  NOR2BX1 U1211 ( .AN(n49), .B(n21), .Y(n523) );
  XNOR2X1 U1212 ( .A(n1), .B(n725), .Y(n707) );
  XNOR2X1 U1213 ( .A(n1), .B(n722), .Y(n709) );
  XNOR2X1 U1214 ( .A(n7), .B(b_10_), .Y(n691) );
  XNOR2X1 U1215 ( .A(n1), .B(n722), .Y(n704) );
  XNOR2X1 U1216 ( .A(n1), .B(n729), .Y(n711) );
  XNOR2X1 U1217 ( .A(b_9_), .B(n1), .Y(n716) );
  XNOR2X1 U1218 ( .A(n728), .B(n1), .Y(n710) );
  XNOR2X1 U1219 ( .A(n726), .B(n1), .Y(n708) );
  XNOR2X1 U1220 ( .A(n726), .B(n7), .Y(n690) );
  XNOR2X1 U1221 ( .A(n735), .B(n1), .Y(n717) );
  XNOR2X1 U1222 ( .A(n731), .B(n7), .Y(n695) );
  XNOR2X1 U1223 ( .A(n732), .B(n13), .Y(n678) );
  XNOR2X1 U1224 ( .A(n733), .B(n13), .Y(n679) );
  XNOR2X1 U1225 ( .A(n735), .B(n19), .Y(n663) );
  XNOR2X1 U1226 ( .A(n730), .B(n7), .Y(n694) );
  XNOR2X1 U1227 ( .A(n723), .B(n1), .Y(n705) );
  XNOR2X1 U1228 ( .A(n730), .B(n31), .Y(n622) );
  XNOR2X1 U1229 ( .A(n721), .B(n1), .Y(n703) );
  ADDHX1 U1230 ( .A(n439), .B(n558), .CO(n431), .S(n432) );
  CLKINVX1 U1231 ( .A(n7), .Y(n768) );
  OAI22XL U1232 ( .A0(n17), .A1(n670), .B0(n669), .B1(n16), .Y(n527) );
  OAI22XL U1233 ( .A0(n699), .A1(n9), .B0(n11), .B1(n700), .Y(n557) );
  OAI22XL U1234 ( .A0(n716), .A1(n5), .B0(n715), .B1(n3), .Y(n573) );
  ADDHXL U1235 ( .A(n564), .B(n548), .CO(n381), .S(n382) );
  OAI22XL U1236 ( .A0(n5), .A1(n707), .B0(n706), .B1(n3), .Y(n564) );
  OAI22XL U1237 ( .A0(n690), .A1(n10), .B0(n12), .B1(n691), .Y(n548) );
  ADDHXL U1238 ( .A(n497), .B(n545), .CO(n351), .S(n352) );
  OAI22XL U1239 ( .A0(n12), .A1(n688), .B0(n687), .B1(n10), .Y(n545) );
  OAI22XL U1240 ( .A0(n29), .A1(n640), .B0(n639), .B1(n27), .Y(n497) );
  ADDHXL U1241 ( .A(n546), .B(n562), .CO(n362), .S(n363) );
  OAI22XL U1242 ( .A0(n5), .A1(n705), .B0(n704), .B1(n3), .Y(n562) );
  OAI22XL U1243 ( .A0(n12), .A1(n689), .B0(n688), .B1(n10), .Y(n546) );
  CLKINVX1 U1244 ( .A(n25), .Y(n765) );
  ADDHXL U1245 ( .A(n438), .B(n540), .CO(n427), .S(n428) );
  OAI22XL U1246 ( .A0(n684), .A1(n16), .B0(n751), .B1(n767), .Y(n438) );
  CLKINVX1 U1247 ( .A(n13), .Y(n767) );
  OAI22XL U1248 ( .A0(n666), .A1(n22), .B0(n24), .B1(n766), .Y(n437) );
  OAI22XL U1249 ( .A0(n713), .A1(n5), .B0(n712), .B1(n3), .Y(n570) );
  CLKINVX1 U1250 ( .A(n19), .Y(n766) );
  CMPR42X1 U1251 ( .A(n530), .B(n363), .C(n370), .D(n498), .ICI(n454), .S(n361), .ICO(n359), .CO(n360) );
  OAI22XL U1252 ( .A0(n593), .A1(n48), .B0(n46), .B1(n592), .Y(n454) );
  OAI22XL U1253 ( .A0(n672), .A1(n16), .B0(n17), .B1(n673), .Y(n530) );
  OAI22XL U1254 ( .A0(n641), .A1(n29), .B0(n640), .B1(n27), .Y(n498) );
  CMPR42X1 U1255 ( .A(n515), .B(n563), .C(n547), .D(n381), .ICI(n499), .S(n372), .ICO(n370), .CO(n371) );
  OAI22XL U1256 ( .A0(n642), .A1(n29), .B0(n641), .B1(n27), .Y(n499) );
  OAI22XL U1257 ( .A0(n753), .A1(n706), .B0(n705), .B1(n3), .Y(n563) );
  OAI22XL U1258 ( .A0(n24), .A1(n658), .B0(n657), .B1(n21), .Y(n515) );
  CMPR42X1 U1259 ( .A(n551), .B(n487), .C(n503), .D(n535), .ICI(n410), .S(n404), .ICO(n402), .CO(n403) );
  OAI22XL U1260 ( .A0(n645), .A1(n27), .B0(n29), .B1(n646), .Y(n503) );
  CMPR42X1 U1261 ( .A(n435), .B(n486), .C(n398), .D(n502), .ICI(n402), .S(n396), .ICO(n394), .CO(n395) );
  OAI22XL U1262 ( .A0(n638), .A1(n27), .B0(n645), .B1(n29), .Y(n502) );
  CMPR42X1 U1263 ( .A(n485), .B(n517), .C(n397), .D(n501), .ICI(n394), .S(n388), .ICO(n386), .CO(n387) );
  OAI22XL U1264 ( .A0(n660), .A1(n24), .B0(n659), .B1(n21), .Y(n517) );
  OAI22XL U1265 ( .A0(n638), .A1(n29), .B0(n643), .B1(n27), .Y(n501) );
  OAI22XL U1266 ( .A0(n627), .A1(n33), .B0(n35), .B1(n628), .Y(n485) );
  CMPR42X1 U1267 ( .A(n500), .B(n470), .C(n389), .D(n484), .ICI(n386), .S(n378), .ICO(n376), .CO(n377) );
  OAI22XL U1268 ( .A0(n611), .A1(n747), .B0(n610), .B1(n40), .Y(n470) );
  OAI22XL U1269 ( .A0(n626), .A1(n33), .B0(n627), .B1(n35), .Y(n484) );
  OAI22XL U1270 ( .A0(n643), .A1(n29), .B0(n642), .B1(n27), .Y(n500) );
  CMPR42X1 U1271 ( .A(n455), .B(n469), .C(n483), .D(n531), .ICI(n376), .S(n369), .ICO(n367), .CO(n368) );
  NOR2BX1 U1272 ( .AN(n49), .B(n46), .Y(n455) );
  OAI22XL U1273 ( .A0(n609), .A1(n40), .B0(n747), .B1(n610), .Y(n469) );
  OAI22XL U1274 ( .A0(n674), .A1(n17), .B0(n673), .B1(n16), .Y(n531) );
  CMPR42X1 U1275 ( .A(n529), .B(n352), .C(n362), .D(n453), .ICI(n359), .S(n350), .ICO(n348), .CO(n349) );
  OAI22XL U1276 ( .A0(n672), .A1(n17), .B0(n671), .B1(n16), .Y(n529) );
  OAI22XL U1277 ( .A0(n591), .A1(n46), .B0(n48), .B1(n592), .Y(n453) );
  CLKBUFX3 U1278 ( .A(n754), .Y(n46) );
  CLKBUFX3 U1279 ( .A(n759), .Y(n16) );
  CLKBUFX3 U1280 ( .A(n853), .Y(n28) );
  CLKBUFX3 U1281 ( .A(n755), .Y(n40) );
  CLKBUFX3 U1282 ( .A(n756), .Y(n34) );
  CLKBUFX3 U1283 ( .A(n760), .Y(n10) );
  CLKBUFX3 U1284 ( .A(n759), .Y(n15) );
  CLKBUFX3 U1285 ( .A(n853), .Y(n27) );
  CLKBUFX3 U1286 ( .A(n756), .Y(n33) );
  CLKBUFX3 U1287 ( .A(n760), .Y(n9) );
  ADDFXL U1288 ( .A(n509), .B(n493), .CI(n310), .CO(n307), .S(n308) );
  OAI22XL U1289 ( .A0(n24), .A1(n652), .B0(n651), .B1(n22), .Y(n509) );
  OAI22XL U1290 ( .A0(n636), .A1(n29), .B0(n635), .B1(n28), .Y(n493) );
  CLKINVX1 U1291 ( .A(n309), .Y(n310) );
  OAI22XL U1292 ( .A0(n659), .A1(n24), .B0(n658), .B1(n21), .Y(n516) );
  CLKINVX1 U1293 ( .A(n37), .Y(n763) );
  CLKBUFX3 U1294 ( .A(n752), .Y(n11) );
  CLKBUFX3 U1295 ( .A(n748), .Y(n35) );
  CLKBUFX3 U1296 ( .A(n761), .Y(n3) );
  CLKBUFX3 U1297 ( .A(n752), .Y(n12) );
  CLKBUFX3 U1298 ( .A(n748), .Y(n36) );
  ADDFXL U1299 ( .A(n569), .B(n505), .CI(n521), .CO(n415), .S(n416) );
  OAI22XL U1300 ( .A0(n5), .A1(n712), .B0(n711), .B1(n3), .Y(n569) );
  OAI22XL U1301 ( .A0(n663), .A1(n21), .B0(n24), .B1(n664), .Y(n521) );
  NOR2BX1 U1302 ( .AN(n49), .B(n27), .Y(n505) );
  OAI22XL U1303 ( .A0(n679), .A1(n17), .B0(n678), .B1(n15), .Y(n536) );
  OAI22XL U1304 ( .A0(n647), .A1(n29), .B0(n646), .B1(n27), .Y(n504) );
  XNOR2X1 U1305 ( .A(n49), .B(n25), .Y(n647) );
  CLKINVX1 U1306 ( .A(n31), .Y(n764) );
  OAI22XL U1307 ( .A0(n24), .A1(n653), .B0(n652), .B1(n22), .Y(n510) );
  CMPR42X1 U1308 ( .A(n291), .B(n475), .C(n490), .D(n461), .ICI(n288), .S(n284), .ICO(n282), .CO(n283) );
  OAI22XL U1309 ( .A0(n600), .A1(n40), .B0(n42), .B1(n601), .Y(n461) );
  OAI22XL U1310 ( .A0(n29), .A1(n633), .B0(n632), .B1(n28), .Y(n490) );
  OAI22XL U1311 ( .A0(n36), .A1(n617), .B0(n616), .B1(n34), .Y(n475) );
  CMPR42X1 U1312 ( .A(n491), .B(n292), .C(n476), .D(n299), .ICI(n296), .S(n290), .ICO(n288), .CO(n289) );
  OAI22XL U1313 ( .A0(n618), .A1(n36), .B0(n617), .B1(n34), .Y(n476) );
  OAI22XL U1314 ( .A0(n29), .A1(n634), .B0(n633), .B1(n28), .Y(n491) );
  CLKINVX1 U1315 ( .A(n291), .Y(n292) );
  ADDFXL U1316 ( .A(n474), .B(n459), .CI(n277), .CO(n270), .S(n271) );
  OAI22XL U1317 ( .A0(n36), .A1(n615), .B0(n614), .B1(n34), .Y(n474) );
  OAI22XL U1318 ( .A0(n42), .A1(n599), .B0(n598), .B1(n40), .Y(n459) );
  ADDFXL U1319 ( .A(n309), .B(n492), .CI(n508), .CO(n299), .S(n300) );
  OAI22XL U1320 ( .A0(n24), .A1(n651), .B0(n650), .B1(n22), .Y(n508) );
  OAI22XL U1321 ( .A0(n29), .A1(n635), .B0(n634), .B1(n28), .Y(n492) );
  CMPR42X1 U1322 ( .A(n443), .B(n458), .C(n265), .D(n262), .ICI(n472), .S(n261), .ICO(n259), .CO(n260) );
  OAI22XL U1323 ( .A0(n42), .A1(n597), .B0(n596), .B1(n40), .Y(n458) );
  OAI22XL U1324 ( .A0(n48), .A1(n581), .B0(n46), .B1(n580), .Y(n443) );
  XNOR2X2 U1325 ( .A(a_5_), .B(a_6_), .Y(n758) );
  XNOR2X1 U1326 ( .A(n1), .B(n724), .Y(n706) );
  XNOR2X1 U1327 ( .A(n1), .B(b_1_), .Y(n718) );
  XNOR2X1 U1328 ( .A(n7), .B(b_1_), .Y(n700) );
  XNOR2X1 U1329 ( .A(n25), .B(b_1_), .Y(n646) );
  XNOR2X1 U1330 ( .A(n19), .B(b_1_), .Y(n664) );
  XNOR2X1 U1331 ( .A(n13), .B(b_1_), .Y(n682) );
  XNOR2X1 U1332 ( .A(n31), .B(b_1_), .Y(n628) );
  XNOR2X1 U1333 ( .A(n37), .B(b_1_), .Y(n610) );
  NAND2X1 U1334 ( .A(n743), .B(n759), .Y(n751) );
  XOR2X1 U1335 ( .A(a_5_), .B(a_4_), .Y(n743) );
  NAND2X1 U1336 ( .A(n742), .B(n758), .Y(n750) );
  XOR2X1 U1337 ( .A(a_7_), .B(a_6_), .Y(n742) );
  NAND2X1 U1338 ( .A(n741), .B(n853), .Y(n749) );
  XOR2X1 U1339 ( .A(a_9_), .B(a_8_), .Y(n741) );
  XOR2X1 U1340 ( .A(a_11_), .B(a_10_), .Y(n740) );
  NAND2X1 U1341 ( .A(n739), .B(n755), .Y(n747) );
  XOR2X1 U1342 ( .A(a_13_), .B(a_12_), .Y(n739) );
  XOR2X1 U1343 ( .A(a_3_), .B(a_2_), .Y(n744) );
  XOR2X1 U1344 ( .A(a_14_), .B(a_15_), .Y(n738) );
  NAND2X1 U1345 ( .A(n745), .B(n761), .Y(n753) );
  XOR2X1 U1346 ( .A(a_0_), .B(a_1_), .Y(n745) );
  XNOR2X1 U1347 ( .A(n31), .B(n724), .Y(n616) );
  XNOR2X1 U1348 ( .A(n43), .B(b_1_), .Y(n592) );
  XNOR2X1 U1349 ( .A(n37), .B(n724), .Y(n598) );
endmodule


module FFT_ultrafast2_shift_DW01_sub_26 ( A, B, DIFF_31_, DIFF_30_, DIFF_29_, 
        DIFF_28_, DIFF_27_, DIFF_26_, DIFF_25_, DIFF_24_, DIFF_23_, DIFF_22_, 
        DIFF_21_, DIFF_20_, DIFF_19_, DIFF_18_, DIFF_17_, DIFF_16_ );
  input [31:0] A;
  input [31:0] B;
  output DIFF_31_, DIFF_30_, DIFF_29_, DIFF_28_, DIFF_27_, DIFF_26_, DIFF_25_,
         DIFF_24_, DIFF_23_, DIFF_22_, DIFF_21_, DIFF_20_, DIFF_19_, DIFF_18_,
         DIFF_17_, DIFF_16_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n19, n22, n24, n25, n26, n27, n28, n30, n32, n33, n34, n35, n36,
         n38, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n54, n56,
         n57, n58, n59, n60, n62, n64, n65, n66, n67, n68, n70, n72, n73, n74,
         n75, n77, n79, n80, n82, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n122, n125, n126, n128, n129, n130, n133, n134, n136, n137,
         n138, n141, n142, n144, n145, n146, n149, n150, n151, n154, n156,
         n158, n160, n162, n164, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308;

  XOR2XL U219 ( .A(n36), .B(n6), .Y(DIFF_27_) );
  OAI21X4 U220 ( .A0(n36), .A1(n34), .B0(n35), .Y(n33) );
  AOI21X4 U221 ( .A0(n41), .A1(n290), .B0(n38), .Y(n36) );
  CLKINVX1 U222 ( .A(B[11]), .Y(n188) );
  OR2X1 U223 ( .A(A[9]), .B(n190), .Y(n307) );
  CLKINVX1 U224 ( .A(B[13]), .Y(n186) );
  CLKINVX1 U225 ( .A(B[15]), .Y(n184) );
  NOR2X1 U226 ( .A(n185), .B(A[14]), .Y(n91) );
  CLKINVX1 U227 ( .A(B[17]), .Y(n182) );
  NAND2X1 U228 ( .A(A[28]), .B(n171), .Y(n32) );
  INVX1 U229 ( .A(n84), .Y(n82) );
  OR2X1 U230 ( .A(n183), .B(A[16]), .Y(n288) );
  NAND2X1 U231 ( .A(n287), .B(n24), .Y(n3) );
  OR2X1 U232 ( .A(n182), .B(A[17]), .Y(n286) );
  OR2X1 U233 ( .A(A[30]), .B(n169), .Y(n287) );
  OR2X1 U234 ( .A(A[28]), .B(n171), .Y(n289) );
  OR2X1 U235 ( .A(A[26]), .B(n173), .Y(n290) );
  OR2X1 U236 ( .A(A[18]), .B(n181), .Y(n291) );
  OR2X1 U237 ( .A(A[20]), .B(n179), .Y(n292) );
  OR2X1 U238 ( .A(A[22]), .B(n177), .Y(n293) );
  OR2X1 U239 ( .A(A[24]), .B(n175), .Y(n294) );
  AND2X2 U240 ( .A(A[9]), .B(n190), .Y(n295) );
  AND2X2 U241 ( .A(n187), .B(A[12]), .Y(n296) );
  AND2X2 U242 ( .A(A[13]), .B(n186), .Y(n297) );
  AND2X2 U243 ( .A(n191), .B(A[8]), .Y(n298) );
  OR2X2 U244 ( .A(n28), .B(n26), .Y(n299) );
  NAND2X2 U245 ( .A(n299), .B(n27), .Y(n25) );
  NAND2X1 U246 ( .A(A[26]), .B(n173), .Y(n40) );
  NOR2X1 U247 ( .A(n170), .B(A[29]), .Y(n26) );
  OR2X1 U248 ( .A(n187), .B(A[12]), .Y(n302) );
  XNOR2X1 U249 ( .A(n25), .B(n3), .Y(DIFF_30_) );
  AOI21X1 U250 ( .A0(n305), .A1(n296), .B0(n297), .Y(n95) );
  AOI21X1 U251 ( .A0(n307), .A1(n298), .B0(n295), .Y(n113) );
  AOI21X4 U252 ( .A0(n33), .A1(n289), .B0(n30), .Y(n28) );
  NAND2X2 U253 ( .A(n170), .B(A[29]), .Y(n27) );
  AO21X4 U254 ( .A0(n25), .A1(n287), .B0(n22), .Y(n300) );
  OAI21X2 U255 ( .A0(n44), .A1(n42), .B0(n43), .Y(n41) );
  OAI21X1 U256 ( .A0(n89), .A1(n92), .B0(n90), .Y(n88) );
  NOR2X1 U257 ( .A(n89), .B(n91), .Y(n87) );
  NOR2XL U258 ( .A(n189), .B(A[10]), .Y(n109) );
  NAND2XL U259 ( .A(n192), .B(A[7]), .Y(n126) );
  NAND2XL U260 ( .A(n195), .B(A[4]), .Y(n137) );
  OAI21X1 U261 ( .A0(n60), .A1(n58), .B0(n59), .Y(n57) );
  OAI21X1 U262 ( .A0(n68), .A1(n66), .B0(n67), .Y(n65) );
  NAND2X1 U263 ( .A(A[30]), .B(n169), .Y(n24) );
  OA21XL U264 ( .A0(n303), .A1(n133), .B0(n134), .Y(n130) );
  OA21XL U265 ( .A0(n138), .A1(n136), .B0(n137), .Y(n303) );
  NAND2XL U266 ( .A(n172), .B(A[27]), .Y(n35) );
  OR2X1 U267 ( .A(n168), .B(A[31]), .Y(n308) );
  OA21XL U268 ( .A0(n306), .A1(n141), .B0(n142), .Y(n138) );
  OA21XL U269 ( .A0(n146), .A1(n144), .B0(n145), .Y(n306) );
  OAI21X2 U270 ( .A0(n52), .A1(n50), .B0(n51), .Y(n49) );
  OAI21X2 U271 ( .A0(n86), .A1(n74), .B0(n75), .Y(n73) );
  XNOR2XL U272 ( .A(n49), .B(n9), .Y(DIFF_24_) );
  NAND2XL U273 ( .A(n294), .B(n48), .Y(n9) );
  XOR2XL U274 ( .A(n52), .B(n10), .Y(DIFF_23_) );
  NAND2XL U275 ( .A(n160), .B(n51), .Y(n10) );
  XNOR2XL U276 ( .A(n57), .B(n11), .Y(DIFF_22_) );
  NAND2XL U277 ( .A(n293), .B(n56), .Y(n11) );
  XOR2XL U278 ( .A(n60), .B(n12), .Y(DIFF_21_) );
  NAND2XL U279 ( .A(n162), .B(n59), .Y(n12) );
  XNOR2XL U280 ( .A(n65), .B(n13), .Y(DIFF_20_) );
  NAND2XL U281 ( .A(n292), .B(n64), .Y(n13) );
  XOR2XL U282 ( .A(n68), .B(n14), .Y(DIFF_19_) );
  NAND2XL U283 ( .A(n164), .B(n67), .Y(n14) );
  XNOR2XL U284 ( .A(n73), .B(n15), .Y(DIFF_18_) );
  NAND2XL U285 ( .A(n291), .B(n72), .Y(n15) );
  NAND2XL U286 ( .A(n286), .B(n79), .Y(n16) );
  AOI21XL U287 ( .A0(n85), .A1(n288), .B0(n82), .Y(n80) );
  NAND2XL U288 ( .A(n288), .B(n84), .Y(n17) );
  INVXL U289 ( .A(n86), .Y(n85) );
  OAI21X1 U290 ( .A0(n104), .A1(n94), .B0(n95), .Y(n93) );
  XNOR2X1 U291 ( .A(n300), .B(n2), .Y(DIFF_31_) );
  NOR2X1 U292 ( .A(n178), .B(A[21]), .Y(n58) );
  NOR2X1 U293 ( .A(n176), .B(A[23]), .Y(n50) );
  NOR2X1 U294 ( .A(n174), .B(A[25]), .Y(n42) );
  NOR2X1 U295 ( .A(n180), .B(A[19]), .Y(n66) );
  NAND2XL U296 ( .A(n184), .B(A[15]), .Y(n90) );
  OR2X1 U297 ( .A(n191), .B(A[8]), .Y(n301) );
  NOR2X1 U298 ( .A(n172), .B(A[27]), .Y(n34) );
  INVX3 U299 ( .A(B[30]), .Y(n169) );
  NAND2XL U300 ( .A(n188), .B(A[11]), .Y(n108) );
  NAND2XL U301 ( .A(n194), .B(A[5]), .Y(n134) );
  NAND2XL U302 ( .A(n196), .B(A[3]), .Y(n142) );
  NAND2XL U303 ( .A(n193), .B(A[6]), .Y(n129) );
  NAND2XL U304 ( .A(A[2]), .B(n197), .Y(n145) );
  NAND2XL U305 ( .A(n198), .B(A[1]), .Y(n150) );
  NOR2BX1 U306 ( .AN(B[0]), .B(A[0]), .Y(n151) );
  AOI21X1 U307 ( .A0(n73), .A1(n291), .B0(n70), .Y(n68) );
  CLKINVX1 U308 ( .A(n72), .Y(n70) );
  AOI21X1 U309 ( .A0(n65), .A1(n292), .B0(n62), .Y(n60) );
  CLKINVX1 U310 ( .A(n64), .Y(n62) );
  AOI21X1 U311 ( .A0(n57), .A1(n293), .B0(n54), .Y(n52) );
  CLKINVX1 U312 ( .A(n56), .Y(n54) );
  AOI21X1 U313 ( .A0(n49), .A1(n294), .B0(n46), .Y(n44) );
  CLKINVX1 U314 ( .A(n48), .Y(n46) );
  CLKINVX1 U315 ( .A(n40), .Y(n38) );
  NAND2X1 U316 ( .A(n288), .B(n286), .Y(n74) );
  AOI21X1 U317 ( .A0(n286), .A1(n82), .B0(n77), .Y(n75) );
  XNOR2X1 U318 ( .A(n41), .B(n7), .Y(DIFF_26_) );
  NAND2X1 U319 ( .A(n290), .B(n40), .Y(n7) );
  XOR2X1 U320 ( .A(n28), .B(n4), .Y(DIFF_29_) );
  NAND2X1 U321 ( .A(n154), .B(n27), .Y(n4) );
  CLKINVX1 U322 ( .A(n26), .Y(n154) );
  XOR2X1 U323 ( .A(n44), .B(n8), .Y(DIFF_25_) );
  NAND2X1 U324 ( .A(n158), .B(n43), .Y(n8) );
  CLKINVX1 U325 ( .A(n42), .Y(n158) );
  CLKINVX1 U326 ( .A(n50), .Y(n160) );
  CLKINVX1 U327 ( .A(n79), .Y(n77) );
  CLKINVX1 U328 ( .A(n24), .Y(n22) );
  CLKINVX1 U329 ( .A(n58), .Y(n162) );
  CLKINVX1 U330 ( .A(n66), .Y(n164) );
  XOR2X1 U331 ( .A(n80), .B(n16), .Y(DIFF_17_) );
  XNOR2X1 U332 ( .A(n85), .B(n17), .Y(DIFF_16_) );
  AOI21X1 U333 ( .A0(n93), .A1(n87), .B0(n88), .Y(n86) );
  CLKINVX1 U334 ( .A(n32), .Y(n30) );
  AOI21X1 U335 ( .A0(n105), .A1(n111), .B0(n106), .Y(n104) );
  OAI21XL U336 ( .A0(n112), .A1(n122), .B0(n113), .Y(n111) );
  NOR2X1 U337 ( .A(n107), .B(n109), .Y(n105) );
  OAI21XL U338 ( .A0(n107), .A1(n110), .B0(n108), .Y(n106) );
  OA21XL U339 ( .A0(n304), .A1(n125), .B0(n126), .Y(n122) );
  OA21XL U340 ( .A0(n130), .A1(n128), .B0(n129), .Y(n304) );
  NOR2X1 U341 ( .A(n184), .B(A[15]), .Y(n89) );
  XNOR2X1 U342 ( .A(n33), .B(n5), .Y(DIFF_28_) );
  NAND2X1 U343 ( .A(n289), .B(n32), .Y(n5) );
  NAND2X1 U344 ( .A(n156), .B(n35), .Y(n6) );
  CLKINVX1 U345 ( .A(n34), .Y(n156) );
  NAND2X1 U346 ( .A(n308), .B(n19), .Y(n2) );
  NAND2X1 U347 ( .A(n182), .B(A[17]), .Y(n79) );
  NAND2X1 U348 ( .A(n183), .B(A[16]), .Y(n84) );
  NAND2X1 U349 ( .A(A[24]), .B(n175), .Y(n48) );
  NAND2X1 U350 ( .A(A[22]), .B(n177), .Y(n56) );
  NAND2X1 U351 ( .A(A[20]), .B(n179), .Y(n64) );
  NAND2X1 U352 ( .A(A[18]), .B(n181), .Y(n72) );
  NAND2X1 U353 ( .A(n174), .B(A[25]), .Y(n43) );
  NAND2X1 U354 ( .A(n176), .B(A[23]), .Y(n51) );
  NAND2X1 U355 ( .A(n178), .B(A[21]), .Y(n59) );
  NAND2X1 U356 ( .A(n180), .B(A[19]), .Y(n67) );
  OR2X1 U357 ( .A(A[13]), .B(n186), .Y(n305) );
  NAND2X1 U358 ( .A(n185), .B(A[14]), .Y(n92) );
  CLKINVX1 U359 ( .A(B[10]), .Y(n189) );
  NOR2X1 U360 ( .A(n188), .B(A[11]), .Y(n107) );
  NOR2X1 U361 ( .A(n192), .B(A[7]), .Y(n125) );
  NOR2X1 U362 ( .A(A[2]), .B(n197), .Y(n144) );
  NOR2X1 U363 ( .A(n196), .B(A[3]), .Y(n141) );
  NOR2X1 U364 ( .A(n194), .B(A[5]), .Y(n133) );
  NOR2X1 U365 ( .A(n195), .B(A[4]), .Y(n136) );
  NAND2X1 U366 ( .A(n168), .B(A[31]), .Y(n19) );
  NOR2X1 U367 ( .A(n193), .B(A[6]), .Y(n128) );
  CLKINVX1 U368 ( .A(B[14]), .Y(n185) );
  CLKINVX1 U369 ( .A(B[26]), .Y(n173) );
  CLKINVX1 U370 ( .A(B[24]), .Y(n175) );
  CLKINVX1 U371 ( .A(B[22]), .Y(n177) );
  CLKINVX1 U372 ( .A(B[20]), .Y(n179) );
  CLKINVX1 U373 ( .A(B[18]), .Y(n181) );
  NAND2X1 U374 ( .A(n189), .B(A[10]), .Y(n110) );
  NAND2X1 U375 ( .A(n307), .B(n301), .Y(n112) );
  NAND2X1 U376 ( .A(n305), .B(n302), .Y(n94) );
  CLKINVX1 U377 ( .A(B[12]), .Y(n187) );
  CLKINVX1 U378 ( .A(B[31]), .Y(n168) );
  CLKINVX1 U379 ( .A(B[16]), .Y(n183) );
  CLKINVX1 U380 ( .A(B[29]), .Y(n170) );
  CLKINVX1 U381 ( .A(B[25]), .Y(n174) );
  CLKINVX1 U382 ( .A(B[23]), .Y(n176) );
  CLKINVX1 U383 ( .A(B[21]), .Y(n178) );
  CLKINVX1 U384 ( .A(B[19]), .Y(n180) );
  CLKINVX1 U385 ( .A(B[3]), .Y(n196) );
  OA21XL U386 ( .A0(n149), .A1(n151), .B0(n150), .Y(n146) );
  CLKINVX1 U387 ( .A(B[1]), .Y(n198) );
  CLKINVX1 U388 ( .A(B[4]), .Y(n195) );
  CLKINVX1 U389 ( .A(B[2]), .Y(n197) );
  NOR2X1 U390 ( .A(n198), .B(A[1]), .Y(n149) );
  CLKINVX1 U391 ( .A(B[6]), .Y(n193) );
  CLKINVX1 U392 ( .A(B[9]), .Y(n190) );
  CLKINVX1 U393 ( .A(B[28]), .Y(n171) );
  CLKINVX1 U394 ( .A(B[5]), .Y(n194) );
  CLKINVX1 U395 ( .A(B[8]), .Y(n191) );
  CLKINVX1 U396 ( .A(B[7]), .Y(n192) );
  CLKINVX1 U397 ( .A(B[27]), .Y(n172) );
endmodule


module FFT_ultrafast2_shift ( clk, rst, fir_valid, fir_d, fft_valid, fft_d1, 
        fft_d2, fft_d3, fft_d4, fft_d5, fft_d6, fft_d7, fft_d8, fft_d9, 
        fft_d10, fft_d11, fft_d12, fft_d13, fft_d14, fft_d15, fft_d0 );
  input [15:0] fir_d;
  output [31:0] fft_d1;
  output [31:0] fft_d2;
  output [31:0] fft_d3;
  output [31:0] fft_d4;
  output [31:0] fft_d5;
  output [31:0] fft_d6;
  output [31:0] fft_d7;
  output [31:0] fft_d8;
  output [31:0] fft_d9;
  output [31:0] fft_d10;
  output [31:0] fft_d11;
  output [31:0] fft_d12;
  output [31:0] fft_d13;
  output [31:0] fft_d14;
  output [31:0] fft_d15;
  output [31:0] fft_d0;
  input clk, rst, fir_valid;
  output fft_valid;
  wire   n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, mul_0_Wn_19, mul_0_Wn_8, mul_0_Wn_6,
         mul_0_Wn_2, mul_0_Wn_1, mul_0_Wn_0, mul_2_Wn_19, mul_2_Wn_11,
         mul_2_Wn_9, mul_2_Wn_8, data_0__15_, data_0__14_, data_0__13_,
         data_0__12_, data_0__11_, data_0__10_, data_0__9_, data_0__8_,
         data_0__7_, data_0__6_, data_0__5_, data_0__4_, data_0__3_,
         data_0__2_, data_0__1_, data_0__0_, data_1__15_, data_1__14_,
         data_1__13_, data_1__12_, data_1__11_, data_1__10_, data_1__9_,
         data_1__8_, data_1__7_, data_1__6_, data_1__5_, data_1__4_,
         data_1__3_, data_1__2_, data_1__1_, data_1__0_, data_2__15_,
         data_2__14_, data_2__13_, data_2__12_, data_2__11_, data_2__10_,
         data_2__9_, data_2__8_, data_2__7_, data_2__6_, data_2__5_,
         data_2__4_, data_2__3_, data_2__2_, data_2__1_, data_2__0_,
         data_3__15_, data_3__14_, data_3__13_, data_3__12_, data_3__11_,
         data_3__10_, data_3__9_, data_3__8_, data_3__7_, data_3__6_,
         data_3__5_, data_3__4_, data_3__3_, data_3__2_, data_3__1_,
         data_3__0_, data_4__15_, data_4__14_, data_4__13_, data_4__12_,
         data_4__11_, data_4__10_, data_4__9_, data_4__8_, data_4__7_,
         data_4__6_, data_4__5_, data_4__4_, data_4__3_, data_4__2_,
         data_4__1_, data_4__0_, data_5__15_, data_5__14_, data_5__13_,
         data_5__12_, data_5__11_, data_5__10_, data_5__9_, data_5__8_,
         data_5__7_, data_5__6_, data_5__5_, data_5__4_, data_5__3_,
         data_5__2_, data_5__1_, data_5__0_, data_6__15_, data_6__14_,
         data_6__13_, data_6__12_, data_6__11_, data_6__10_, data_6__9_,
         data_6__8_, data_6__7_, data_6__6_, data_6__5_, data_6__4_,
         data_6__3_, data_6__2_, data_6__1_, data_6__0_, data_7__15_,
         data_7__14_, data_7__13_, data_7__12_, data_7__11_, data_7__10_,
         data_7__9_, data_7__8_, data_7__7_, data_7__6_, data_7__5_,
         data_7__4_, data_7__3_, data_7__2_, data_7__1_, data_7__0_,
         data_8__15_, data_8__14_, data_8__13_, data_8__12_, data_8__11_,
         data_8__10_, data_8__9_, data_8__8_, data_8__7_, data_8__6_,
         data_8__5_, data_8__4_, data_8__3_, data_8__2_, data_8__1_,
         data_8__0_, data_9__15_, data_9__14_, data_9__13_, data_9__12_,
         data_9__11_, data_9__10_, data_9__9_, data_9__8_, data_9__7_,
         data_9__6_, data_9__5_, data_9__4_, data_9__3_, data_9__2_,
         data_9__1_, data_9__0_, data_10__15_, data_10__14_, data_10__13_,
         data_10__12_, data_10__11_, data_10__10_, data_10__9_, data_10__8_,
         data_10__7_, data_10__6_, data_10__5_, data_10__4_, data_10__3_,
         data_10__2_, data_10__1_, data_10__0_, data_11__15_, data_11__14_,
         data_11__13_, data_11__12_, data_11__11_, data_11__10_, data_11__9_,
         data_11__8_, data_11__7_, data_11__6_, data_11__5_, data_11__4_,
         data_11__3_, data_11__2_, data_11__1_, data_11__0_, data_12__15_,
         data_12__14_, data_12__13_, data_12__12_, data_12__11_, data_12__10_,
         data_12__9_, data_12__8_, data_12__7_, data_12__6_, data_12__5_,
         data_12__4_, data_12__3_, data_12__2_, data_12__1_, data_12__0_,
         data_13__15_, data_13__14_, data_13__13_, data_13__12_, data_13__11_,
         data_13__10_, data_13__9_, data_13__8_, data_13__7_, data_13__6_,
         data_13__5_, data_13__4_, data_13__3_, data_13__2_, data_13__1_,
         data_13__0_, data_14__15_, data_14__14_, data_14__13_, data_14__12_,
         data_14__11_, data_14__10_, data_14__9_, data_14__8_, data_14__7_,
         data_14__6_, data_14__5_, data_14__4_, data_14__3_, data_14__2_,
         data_14__1_, data_14__0_, stg1_real_0__15_, stg1_real_0__14_,
         stg1_real_0__13_, stg1_real_0__12_, stg1_real_0__11_,
         stg1_real_0__10_, stg1_real_0__9_, stg1_real_0__8_, stg1_real_0__7_,
         stg1_real_0__6_, stg1_real_0__5_, stg1_real_0__4_, stg1_real_0__3_,
         stg1_real_0__2_, stg1_real_0__1_, stg1_real_0__0_, stg1_real_1__15_,
         stg1_real_1__14_, stg1_real_1__13_, stg1_real_1__12_,
         stg1_real_1__11_, stg1_real_1__10_, stg1_real_1__9_, stg1_real_1__8_,
         stg1_real_1__7_, stg1_real_1__6_, stg1_real_1__5_, stg1_real_1__4_,
         stg1_real_1__3_, stg1_real_1__2_, stg1_real_1__1_, stg1_real_1__0_,
         stg1_real_2__15_, stg1_real_2__14_, stg1_real_2__13_,
         stg1_real_2__12_, stg1_real_2__11_, stg1_real_2__10_, stg1_real_2__9_,
         stg1_real_2__8_, stg1_real_2__7_, stg1_real_2__6_, stg1_real_2__5_,
         stg1_real_2__4_, stg1_real_2__3_, stg1_real_2__2_, stg1_real_2__1_,
         stg1_real_2__0_, stg1_real_3__15_, stg1_real_3__14_, stg1_real_3__13_,
         stg1_real_3__12_, stg1_real_3__11_, stg1_real_3__10_, stg1_real_3__9_,
         stg1_real_3__8_, stg1_real_3__7_, stg1_real_3__6_, stg1_real_3__5_,
         stg1_real_3__4_, stg1_real_3__3_, stg1_real_3__2_, stg1_real_3__1_,
         stg1_real_3__0_, stg1_real_4__15_, stg1_real_4__14_, stg1_real_4__13_,
         stg1_real_4__12_, stg1_real_4__11_, stg1_real_4__10_, stg1_real_4__9_,
         stg1_real_4__8_, stg1_real_4__7_, stg1_real_4__6_, stg1_real_4__5_,
         stg1_real_4__4_, stg1_real_4__3_, stg1_real_4__2_, stg1_real_4__1_,
         stg1_real_4__0_, stg1_real_5__15_, stg1_real_5__14_, stg1_real_5__13_,
         stg1_real_5__12_, stg1_real_5__11_, stg1_real_5__10_, stg1_real_5__9_,
         stg1_real_5__8_, stg1_real_5__7_, stg1_real_5__6_, stg1_real_5__5_,
         stg1_real_5__4_, stg1_real_5__3_, stg1_real_5__2_, stg1_real_5__1_,
         stg1_real_5__0_, stg1_real_6__15_, stg1_real_6__14_, stg1_real_6__13_,
         stg1_real_6__12_, stg1_real_6__11_, stg1_real_6__10_, stg1_real_6__9_,
         stg1_real_6__8_, stg1_real_6__7_, stg1_real_6__6_, stg1_real_6__5_,
         stg1_real_6__4_, stg1_real_6__3_, stg1_real_6__2_, stg1_real_6__1_,
         stg1_real_6__0_, stg1_real_7__15_, stg1_real_7__14_, stg1_real_7__13_,
         stg1_real_7__12_, stg1_real_7__11_, stg1_real_7__10_, stg1_real_7__9_,
         stg1_real_7__8_, stg1_real_7__7_, stg1_real_7__6_, stg1_real_7__5_,
         stg1_real_7__4_, stg1_real_7__3_, stg1_real_7__2_, stg1_real_7__1_,
         stg1_real_7__0_, stg2_real_0__15_, stg2_real_0__14_, stg2_real_0__13_,
         stg2_real_0__12_, stg2_real_0__11_, stg2_real_0__10_, stg2_real_0__9_,
         stg2_real_0__8_, stg2_real_0__7_, stg2_real_0__6_, stg2_real_0__5_,
         stg2_real_0__4_, stg2_real_0__3_, stg2_real_0__2_, stg2_real_0__1_,
         stg2_real_0__0_, stg2_real_1__15_, stg2_real_1__14_, stg2_real_1__13_,
         stg2_real_1__12_, stg2_real_1__11_, stg2_real_1__10_, stg2_real_1__9_,
         stg2_real_1__8_, stg2_real_1__7_, stg2_real_1__6_, stg2_real_1__5_,
         stg2_real_1__4_, stg2_real_1__3_, stg2_real_1__2_, stg2_real_1__1_,
         stg2_real_1__0_, stg2_real_2__15_, stg2_real_2__14_, stg2_real_2__13_,
         stg2_real_2__12_, stg2_real_2__11_, stg2_real_2__10_, stg2_real_2__9_,
         stg2_real_2__8_, stg2_real_2__7_, stg2_real_2__6_, stg2_real_2__5_,
         stg2_real_2__4_, stg2_real_2__3_, stg2_real_2__2_, stg2_real_2__1_,
         stg2_real_2__0_, stg2_real_3__15_, stg2_real_3__14_, stg2_real_3__13_,
         stg2_real_3__12_, stg2_real_3__11_, stg2_real_3__10_, stg2_real_3__9_,
         stg2_real_3__8_, stg2_real_3__7_, stg2_real_3__6_, stg2_real_3__5_,
         stg2_real_3__4_, stg2_real_3__3_, stg2_real_3__2_, stg2_real_3__1_,
         stg2_real_3__0_, stg2_real_4__15_, stg2_real_4__14_, stg2_real_4__13_,
         stg2_real_4__12_, stg2_real_4__11_, stg2_real_4__10_, stg2_real_4__9_,
         stg2_real_4__8_, stg2_real_4__7_, stg2_real_4__6_, stg2_real_4__5_,
         stg2_real_4__4_, stg2_real_4__3_, stg2_real_4__2_, stg2_real_4__1_,
         stg2_real_4__0_, stg2_real_5__15_, stg2_real_5__14_, stg2_real_5__13_,
         stg2_real_5__12_, stg2_real_5__11_, stg2_real_5__10_, stg2_real_5__9_,
         stg2_real_5__8_, stg2_real_5__7_, stg2_real_5__6_, stg2_real_5__5_,
         stg2_real_5__4_, stg2_real_5__3_, stg2_real_5__2_, stg2_real_5__1_,
         stg2_real_5__0_, stg2_real_6__15_, stg2_real_6__14_, stg2_real_6__13_,
         stg2_real_6__12_, stg2_real_6__11_, stg2_real_6__10_, stg2_real_6__9_,
         stg2_real_6__8_, stg2_real_6__7_, stg2_real_6__6_, stg2_real_6__5_,
         stg2_real_6__4_, stg2_real_6__3_, stg2_real_6__2_, stg2_real_6__1_,
         stg2_real_6__0_, stg2_real_7__15_, stg2_real_7__14_, stg2_real_7__13_,
         stg2_real_7__12_, stg2_real_7__11_, stg2_real_7__10_, stg2_real_7__9_,
         stg2_real_7__8_, stg2_real_7__7_, stg2_real_7__6_, stg2_real_7__5_,
         stg2_real_7__4_, stg2_real_7__3_, stg2_real_7__2_, stg2_real_7__1_,
         stg2_real_7__0_, stg2_real_12__15_, stg2_real_12__14_,
         stg2_real_12__13_, stg2_real_12__12_, stg2_real_12__11_,
         stg2_real_12__10_, stg2_real_12__9_, stg2_real_12__8_,
         stg2_real_12__7_, stg2_real_12__6_, stg2_real_12__5_,
         stg2_real_12__4_, stg2_real_12__3_, stg2_real_12__2_,
         stg2_real_12__1_, stg2_real_12__0_, stg2_real_13__15_,
         stg2_real_13__14_, stg2_real_13__13_, stg2_real_13__12_,
         stg2_real_13__11_, stg2_real_13__10_, stg2_real_13__9_,
         stg2_real_13__8_, stg2_real_13__7_, stg2_real_13__6_,
         stg2_real_13__5_, stg2_real_13__4_, stg2_real_13__3_,
         stg2_real_13__2_, stg2_real_13__1_, stg2_real_13__0_,
         stg2_real_14__15_, stg2_real_14__14_, stg2_real_14__13_,
         stg2_real_14__12_, stg2_real_14__11_, stg2_real_14__10_,
         stg2_real_14__9_, stg2_real_14__8_, stg2_real_14__7_,
         stg2_real_14__6_, stg2_real_14__5_, stg2_real_14__4_,
         stg2_real_14__3_, stg2_real_14__2_, stg2_real_14__1_,
         stg2_real_14__0_, stg2_real_15__15_, stg2_real_15__14_,
         stg2_real_15__13_, stg2_real_15__12_, stg2_real_15__11_,
         stg2_real_15__10_, stg2_real_15__9_, stg2_real_15__8_,
         stg2_real_15__7_, stg2_real_15__6_, stg2_real_15__5_,
         stg2_real_15__4_, stg2_real_15__3_, stg2_real_15__2_,
         stg2_real_15__1_, stg2_real_15__0_, stg2_img_8__15_, stg2_img_8__14_,
         stg2_img_8__13_, stg2_img_8__12_, stg2_img_8__11_, stg2_img_8__10_,
         stg2_img_8__9_, stg2_img_8__8_, stg2_img_8__7_, stg2_img_8__6_,
         stg2_img_8__5_, stg2_img_8__4_, stg2_img_8__3_, stg2_img_8__2_,
         stg2_img_8__1_, stg2_img_8__0_, stg2_img_9__15_, stg2_img_9__14_,
         stg2_img_9__13_, stg2_img_9__12_, stg2_img_9__11_, stg2_img_9__10_,
         stg2_img_9__9_, stg2_img_9__8_, stg2_img_9__7_, stg2_img_9__6_,
         stg2_img_9__5_, stg2_img_9__4_, stg2_img_9__3_, stg2_img_9__2_,
         stg2_img_9__1_, stg2_img_10__15_, stg2_img_10__14_, stg2_img_10__13_,
         stg2_img_10__12_, stg2_img_10__11_, stg2_img_10__10_, stg2_img_10__9_,
         stg2_img_10__8_, stg2_img_10__7_, stg2_img_10__6_, stg2_img_10__5_,
         stg2_img_10__4_, stg2_img_10__3_, stg2_img_10__2_, stg2_img_10__1_,
         stg2_img_11__15_, stg2_img_11__14_, stg2_img_11__13_,
         stg2_img_11__12_, stg2_img_11__11_, stg2_img_11__10_, stg2_img_11__9_,
         stg2_img_11__8_, stg2_img_11__7_, stg2_img_11__6_, stg2_img_11__5_,
         stg2_img_11__4_, stg2_img_11__3_, stg2_img_11__2_, stg2_img_11__1_,
         stg2_img_13__15_, stg2_img_13__14_, stg2_img_13__13_,
         stg2_img_13__12_, stg2_img_13__11_, stg2_img_13__10_, stg2_img_13__9_,
         stg2_img_13__8_, stg2_img_13__7_, stg2_img_13__6_, stg2_img_13__5_,
         stg2_img_13__4_, stg2_img_13__3_, stg2_img_13__2_, stg2_img_13__1_,
         stg2_img_13__0_, stg2_img_14__15_, stg2_img_14__14_, stg2_img_14__13_,
         stg2_img_14__12_, stg2_img_14__11_, stg2_img_14__10_, stg2_img_14__9_,
         stg2_img_14__8_, stg2_img_14__7_, stg2_img_14__6_, stg2_img_14__5_,
         stg2_img_14__4_, stg2_img_14__3_, stg2_img_14__2_, stg2_img_14__1_,
         stg2_img_14__0_, stg2_img_15__15_, stg2_img_15__14_, stg2_img_15__13_,
         stg2_img_15__12_, stg2_img_15__11_, stg2_img_15__10_, stg2_img_15__9_,
         stg2_img_15__8_, stg2_img_15__7_, stg2_img_15__6_, stg2_img_15__5_,
         stg2_img_15__4_, stg2_img_15__3_, stg2_img_15__2_, stg2_img_15__1_,
         stg2_img_15__0_, N36, N37, N38, N39, N663, N664, N665, N666, N667,
         N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678,
         N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689,
         N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722,
         N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733,
         N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744,
         N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755,
         N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766,
         N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777,
         N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788,
         N789, N790, N919, N920, N921, N922, N923, N924, N925, N926, N927,
         N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938,
         N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949,
         N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960,
         N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971,
         N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982,
         N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993,
         N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034,
         N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044,
         N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054,
         N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064,
         N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074,
         N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084,
         N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094,
         N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104,
         N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114,
         N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124,
         N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134,
         N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1810, n1811, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, mul_1_out_9_, mul_1_out_8_, mul_1_out_7_, mul_1_out_6_,
         mul_1_out_5_, mul_1_out_4_, mul_1_out_3_, mul_1_out_31_,
         mul_1_out_30_, mul_1_out_2_, mul_1_out_29_, mul_1_out_28_,
         mul_1_out_27_, mul_1_out_26_, mul_1_out_25_, mul_1_out_24_,
         mul_1_out_23_, mul_1_out_22_, mul_1_out_21_, mul_1_out_20_,
         mul_1_out_1_, mul_1_out_19_, mul_1_out_18_, mul_1_out_17_,
         mul_1_out_16_, mul_1_out_15_, mul_1_out_14_, mul_1_out_13_,
         mul_1_out_12_, mul_1_out_11_, mul_1_out_10_, mul_1_out_0_,
         mul_0_out_9_, mul_0_out_8_, mul_0_out_7_, mul_0_out_6_, mul_0_out_5_,
         mul_0_out_4_, mul_0_out_3_, mul_0_out_31_, mul_0_out_30_,
         mul_0_out_2_, mul_0_out_29_, mul_0_out_28_, mul_0_out_27_,
         mul_0_out_26_, mul_0_out_25_, mul_0_out_24_, mul_0_out_23_,
         mul_0_out_22_, mul_0_out_21_, mul_0_out_20_, mul_0_out_1_,
         mul_0_out_19_, mul_0_out_18_, mul_0_out_17_, mul_0_out_16_,
         mul_0_out_15_, mul_0_out_14_, mul_0_out_13_, mul_0_out_12_,
         mul_0_out_11_, mul_0_out_10_, mul_0_out_0_, mul_3_out_9_,
         mul_3_out_8_, mul_3_out_7_, mul_3_out_6_, mul_3_out_5_, mul_3_out_4_,
         mul_3_out_3_, mul_3_out_31_, mul_3_out_30_, mul_3_out_2_,
         mul_3_out_29_, mul_3_out_28_, mul_3_out_27_, mul_3_out_26_,
         mul_3_out_25_, mul_3_out_24_, mul_3_out_23_, mul_3_out_22_,
         mul_3_out_21_, mul_3_out_20_, mul_3_out_1_, mul_3_out_19_,
         mul_3_out_18_, mul_3_out_17_, mul_3_out_16_, mul_3_out_15_,
         mul_3_out_14_, mul_3_out_13_, mul_3_out_12_, mul_3_out_11_,
         mul_3_out_10_, mul_3_out_0_, mul_2_out_9_, mul_2_out_8_, mul_2_out_7_,
         mul_2_out_6_, mul_2_out_5_, mul_2_out_4_, mul_2_out_3_, mul_2_out_31_,
         mul_2_out_30_, mul_2_out_2_, mul_2_out_29_, mul_2_out_28_,
         mul_2_out_27_, mul_2_out_26_, mul_2_out_25_, mul_2_out_24_,
         mul_2_out_23_, mul_2_out_22_, mul_2_out_21_, mul_2_out_20_,
         mul_2_out_1_, mul_2_out_19_, mul_2_out_18_, mul_2_out_17_,
         mul_2_out_16_, mul_2_out_15_, mul_2_out_14_, mul_2_out_13_,
         mul_2_out_12_, mul_2_out_11_, mul_2_out_10_, mul_2_out_0_, n17, n18,
         n19, n20, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n339, n341, n468, n7160, n7200, n7220, n7240, n7250,
         n7260, n7270, n7280, n7290, n7300, n7310, n7320, n7330, n7340, n7350,
         n7360, n7370, n7380, n7390, n7400, n7410, n7420, n7430, n7440, n7450,
         n7460, n7470, n7480, n7490, n7500, n7510, n7520, n7530, n7540, n7550,
         n7560, n7570, n7580, n7590, n7600, n7610, n7620, n7630, n7640, n7650,
         n7660, n7670, n7680, n7690, n7700, n7710, n7720, n7730, n7740, n7750,
         n7760, n7770, n7780, n7790, n7800, n7810, n7820, n7830, n7840, n7850,
         n7860, n7870, n7880, n7890, n7900, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n9190, n9200, n9210, n9220, n9230, n9240, n9250, n9260, n9270,
         n9280, n9290, n9300, n9310, n9320, n9330, n9340, n9350, n9360, n9370,
         n9380, n9390, n9400, n9410, n9420, n9430, n9440, n9450, n9460, n9470,
         n9480, n9490, n9500, n9510, n9520, n9530, n9540, n9550, n9560, n9570,
         n9580, n9590, n9600, n9610, n9620, n9630, n9640, n9650, n9660, n9670,
         n9680, n9690, n9700, n9710, n9720, n9730, n9740, n9750, n9760, n9770,
         n9780, n9790, n9800, n9810, n9820, n9830, n9840, n9850, n9860, n9870,
         n9880, n9890, n9900, n9910, n9920, n9930, n9940, n9950, n9960, n9970,
         n9980, n9990, n10000, n10010, n10020, n10030, n10040, n10050, n10060,
         n10070, n10080, n10090, n10100, n10110, n10120, n10130, n10140,
         n10150, n10160, n10170, n10180, n10190, n10200, n10210, n10220,
         n10230, n10240, n10250, n10260, n10270, n10280, n10290, n10300,
         n10310, n10320, n10330, n10340, n10350, n10360, n10370, n10380,
         n10390, n10400, n10410, n10420, n10430, n10440, n10450, n10460,
         n10470, n10480, n10490, n10500, n10510, n10520, n10530, n10540,
         n10550, n10560, n10570, n10580, n10590, n10600, n10610, n10620,
         n10630, n10640, n10650, n10660, n10670, n10680, n10690, n10700,
         n10710, n10720, n10730, n10740, n10750, n10760, n10770, n10780,
         n10790, n10800, n10810, n10820, n10830, n10840, n10850, n10860,
         n10870, n10880, n10890, n10900, n10910, n10920, n10930, n10940,
         n10950, n10960, n10970, n10980, n10990, n11000, n11010, n11020,
         n11030, n11040, n11050, n11060, n11070, n11080, n11090, n11100,
         n11110, n11120, n11130, n11140, n11150, n11160, n11170, n11180,
         n11190, n11200, n11210, n11220, n11230, n11240, n11250, n11260,
         n11270, n11280, n11290, n11300, n11310, n11320, n11330, n11340,
         n11350, n11360, n11370, n11380, n11390, n11400, n11410, n11420, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1812, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224;
  wire   [15:11] mul_0_Wn;
  wire   [15:0] mul_1_in;
  wire   [31:16] mul_o_sub;
  wire   [15:0] mul_2_in;
  wire   [14:13] mul_2_Wn;
  wire   [31:16] mul_o_add;
  wire   [63:0] stg2_real_Wn;
  wire   [63:0] stg3_real;
  wire   [63:0] stg2_img_Wn;
  wire   [63:0] stg3_img;
  wire   [63:0] stg4_real;
  wire   [63:0] stg4_img;
  wire   [159:0] stg_reg;

  FFT_ultrafast2_shift_DW01_sub_0 sub_387 ( .A(stg3_img[31:16]), .B(
        stg3_img[15:0]), .DIFF(stg4_img[15:0]) );
  FFT_ultrafast2_shift_DW01_add_0 add_386 ( .A(stg3_img[31:16]), .B(
        stg3_img[15:0]), .SUM(stg4_img[31:16]) );
  FFT_ultrafast2_shift_DW01_sub_1 sub_385 ( .A(stg3_img[63:48]), .B(
        stg3_img[47:32]), .DIFF(stg4_img[47:32]) );
  FFT_ultrafast2_shift_DW01_add_1 add_384 ( .A(stg3_img[63:48]), .B(
        stg3_img[47:32]), .SUM(stg4_img[63:48]) );
  FFT_ultrafast2_shift_DW01_sub_2 sub_382 ( .A(stg3_real[31:16]), .B(
        stg3_real[15:0]), .DIFF(stg4_real[15:0]) );
  FFT_ultrafast2_shift_DW01_add_2 add_381 ( .A(stg3_real[31:16]), .B(
        stg3_real[15:0]), .SUM(stg4_real[31:16]) );
  FFT_ultrafast2_shift_DW01_sub_3 sub_380 ( .A(stg3_real[63:48]), .B(
        stg3_real[47:32]), .DIFF(stg4_real[47:32]) );
  FFT_ultrafast2_shift_DW01_add_3 add_379 ( .A(stg3_real[63:48]), .B(
        stg3_real[47:32]), .SUM(stg4_real[63:48]) );
  FFT_ultrafast2_shift_DW01_sub_4 sub_365 ( .A(stg2_real_Wn[15:0]), .B(
        stg2_real_Wn[47:32]), .DIFF(stg3_img[15:0]) );
  FFT_ultrafast2_shift_DW01_sub_5 sub_364 ( .A(stg2_img_Wn[63:48]), .B(
        stg2_img_Wn[31:16]), .DIFF(stg3_img[31:16]) );
  FFT_ultrafast2_shift_DW01_add_4 add_363 ( .A(stg2_img_Wn[47:32]), .B(
        stg2_img_Wn[15:0]), .SUM(stg3_img[47:32]) );
  FFT_ultrafast2_shift_DW01_add_5 add_362 ( .A(stg2_img_Wn[63:48]), .B(
        stg2_img_Wn[31:16]), .SUM(stg3_img[63:48]) );
  FFT_ultrafast2_shift_DW01_sub_6 sub_348 ( .A(stg2_img_Wn[47:32]), .B(
        stg2_img_Wn[15:0]), .DIFF(stg3_real[15:0]) );
  FFT_ultrafast2_shift_DW01_sub_7 sub_347 ( .A(stg2_real_Wn[63:48]), .B(
        stg2_real_Wn[31:16]), .DIFF(stg3_real[31:16]) );
  FFT_ultrafast2_shift_DW01_add_6 add_346 ( .A(stg2_real_Wn[47:32]), .B(
        stg2_real_Wn[15:0]), .SUM(stg3_real[47:32]) );
  FFT_ultrafast2_shift_DW01_add_7 add_345 ( .A(stg2_real_Wn[63:48]), .B(
        stg2_real_Wn[31:16]), .SUM(stg3_real[63:48]) );
  FFT_ultrafast2_shift_DW01_sub_12 sub_317 ( .A({stg1_real_3__15_, 
        stg1_real_3__14_, stg1_real_3__13_, stg1_real_3__12_, stg1_real_3__11_, 
        stg1_real_3__10_, stg1_real_3__9_, stg1_real_3__8_, stg1_real_3__7_, 
        stg1_real_3__6_, stg1_real_3__5_, stg1_real_3__4_, stg1_real_3__3_, 
        stg1_real_3__2_, stg1_real_3__1_, stg1_real_3__0_}), .B({
        stg1_real_7__15_, stg1_real_7__14_, stg1_real_7__13_, stg1_real_7__12_, 
        stg1_real_7__11_, stg1_real_7__10_, stg1_real_7__9_, stg1_real_7__8_, 
        stg1_real_7__7_, stg1_real_7__6_, stg1_real_7__5_, stg1_real_7__4_, 
        stg1_real_7__3_, stg1_real_7__2_, stg1_real_7__1_, stg1_real_7__0_}), 
        .DIFF({stg2_real_7__15_, stg2_real_7__14_, stg2_real_7__13_, 
        stg2_real_7__12_, stg2_real_7__11_, stg2_real_7__10_, stg2_real_7__9_, 
        stg2_real_7__8_, stg2_real_7__7_, stg2_real_7__6_, stg2_real_7__5_, 
        stg2_real_7__4_, stg2_real_7__3_, stg2_real_7__2_, stg2_real_7__1_, 
        stg2_real_7__0_}) );
  FFT_ultrafast2_shift_DW01_sub_13 sub_316 ( .A({stg1_real_2__15_, 
        stg1_real_2__14_, stg1_real_2__13_, stg1_real_2__12_, stg1_real_2__11_, 
        stg1_real_2__10_, stg1_real_2__9_, stg1_real_2__8_, stg1_real_2__7_, 
        stg1_real_2__6_, stg1_real_2__5_, stg1_real_2__4_, stg1_real_2__3_, 
        stg1_real_2__2_, stg1_real_2__1_, stg1_real_2__0_}), .B({
        stg1_real_6__15_, stg1_real_6__14_, stg1_real_6__13_, stg1_real_6__12_, 
        stg1_real_6__11_, stg1_real_6__10_, stg1_real_6__9_, stg1_real_6__8_, 
        stg1_real_6__7_, stg1_real_6__6_, stg1_real_6__5_, stg1_real_6__4_, 
        stg1_real_6__3_, stg1_real_6__2_, stg1_real_6__1_, stg1_real_6__0_}), 
        .DIFF({stg2_real_6__15_, stg2_real_6__14_, stg2_real_6__13_, 
        stg2_real_6__12_, stg2_real_6__11_, stg2_real_6__10_, stg2_real_6__9_, 
        stg2_real_6__8_, stg2_real_6__7_, stg2_real_6__6_, stg2_real_6__5_, 
        stg2_real_6__4_, stg2_real_6__3_, stg2_real_6__2_, stg2_real_6__1_, 
        stg2_real_6__0_}) );
  FFT_ultrafast2_shift_DW01_sub_14 sub_315 ( .A({stg1_real_1__15_, 
        stg1_real_1__14_, stg1_real_1__13_, stg1_real_1__12_, stg1_real_1__11_, 
        stg1_real_1__10_, stg1_real_1__9_, stg1_real_1__8_, stg1_real_1__7_, 
        stg1_real_1__6_, stg1_real_1__5_, stg1_real_1__4_, stg1_real_1__3_, 
        stg1_real_1__2_, stg1_real_1__1_, stg1_real_1__0_}), .B({
        stg1_real_5__15_, stg1_real_5__14_, stg1_real_5__13_, stg1_real_5__12_, 
        stg1_real_5__11_, stg1_real_5__10_, stg1_real_5__9_, stg1_real_5__8_, 
        stg1_real_5__7_, stg1_real_5__6_, stg1_real_5__5_, stg1_real_5__4_, 
        stg1_real_5__3_, stg1_real_5__2_, stg1_real_5__1_, stg1_real_5__0_}), 
        .DIFF({stg2_real_5__15_, stg2_real_5__14_, stg2_real_5__13_, 
        stg2_real_5__12_, stg2_real_5__11_, stg2_real_5__10_, stg2_real_5__9_, 
        stg2_real_5__8_, stg2_real_5__7_, stg2_real_5__6_, stg2_real_5__5_, 
        stg2_real_5__4_, stg2_real_5__3_, stg2_real_5__2_, stg2_real_5__1_, 
        stg2_real_5__0_}) );
  FFT_ultrafast2_shift_DW01_sub_15 sub_314 ( .A({stg1_real_0__15_, 
        stg1_real_0__14_, stg1_real_0__13_, stg1_real_0__12_, stg1_real_0__11_, 
        stg1_real_0__10_, stg1_real_0__9_, stg1_real_0__8_, stg1_real_0__7_, 
        stg1_real_0__6_, stg1_real_0__5_, stg1_real_0__4_, stg1_real_0__3_, 
        stg1_real_0__2_, stg1_real_0__1_, stg1_real_0__0_}), .B({
        stg1_real_4__15_, stg1_real_4__14_, stg1_real_4__13_, stg1_real_4__12_, 
        stg1_real_4__11_, stg1_real_4__10_, stg1_real_4__9_, stg1_real_4__8_, 
        stg1_real_4__7_, stg1_real_4__6_, stg1_real_4__5_, stg1_real_4__4_, 
        stg1_real_4__3_, stg1_real_4__2_, stg1_real_4__1_, stg1_real_4__0_}), 
        .DIFF({stg2_real_4__15_, stg2_real_4__14_, stg2_real_4__13_, 
        stg2_real_4__12_, stg2_real_4__11_, stg2_real_4__10_, stg2_real_4__9_, 
        stg2_real_4__8_, stg2_real_4__7_, stg2_real_4__6_, stg2_real_4__5_, 
        stg2_real_4__4_, stg2_real_4__3_, stg2_real_4__2_, stg2_real_4__1_, 
        stg2_real_4__0_}) );
  FFT_ultrafast2_shift_DW01_add_8 add_313 ( .A({stg1_real_3__15_, 
        stg1_real_3__14_, stg1_real_3__13_, stg1_real_3__12_, stg1_real_3__11_, 
        stg1_real_3__10_, stg1_real_3__9_, stg1_real_3__8_, stg1_real_3__7_, 
        stg1_real_3__6_, stg1_real_3__5_, stg1_real_3__4_, stg1_real_3__3_, 
        stg1_real_3__2_, stg1_real_3__1_, stg1_real_3__0_}), .B({
        stg1_real_7__15_, stg1_real_7__14_, stg1_real_7__13_, stg1_real_7__12_, 
        stg1_real_7__11_, stg1_real_7__10_, stg1_real_7__9_, stg1_real_7__8_, 
        stg1_real_7__7_, stg1_real_7__6_, stg1_real_7__5_, stg1_real_7__4_, 
        stg1_real_7__3_, stg1_real_7__2_, stg1_real_7__1_, stg1_real_7__0_}), 
        .SUM({stg2_real_3__15_, stg2_real_3__14_, stg2_real_3__13_, 
        stg2_real_3__12_, stg2_real_3__11_, stg2_real_3__10_, stg2_real_3__9_, 
        stg2_real_3__8_, stg2_real_3__7_, stg2_real_3__6_, stg2_real_3__5_, 
        stg2_real_3__4_, stg2_real_3__3_, stg2_real_3__2_, stg2_real_3__1_, 
        stg2_real_3__0_}) );
  FFT_ultrafast2_shift_DW01_add_9 add_312 ( .A({stg1_real_2__15_, 
        stg1_real_2__14_, stg1_real_2__13_, stg1_real_2__12_, stg1_real_2__11_, 
        stg1_real_2__10_, stg1_real_2__9_, stg1_real_2__8_, stg1_real_2__7_, 
        stg1_real_2__6_, stg1_real_2__5_, stg1_real_2__4_, stg1_real_2__3_, 
        stg1_real_2__2_, stg1_real_2__1_, stg1_real_2__0_}), .B({
        stg1_real_6__15_, stg1_real_6__14_, stg1_real_6__13_, stg1_real_6__12_, 
        stg1_real_6__11_, stg1_real_6__10_, stg1_real_6__9_, stg1_real_6__8_, 
        stg1_real_6__7_, stg1_real_6__6_, stg1_real_6__5_, stg1_real_6__4_, 
        stg1_real_6__3_, stg1_real_6__2_, stg1_real_6__1_, stg1_real_6__0_}), 
        .SUM({stg2_real_2__15_, stg2_real_2__14_, stg2_real_2__13_, 
        stg2_real_2__12_, stg2_real_2__11_, stg2_real_2__10_, stg2_real_2__9_, 
        stg2_real_2__8_, stg2_real_2__7_, stg2_real_2__6_, stg2_real_2__5_, 
        stg2_real_2__4_, stg2_real_2__3_, stg2_real_2__2_, stg2_real_2__1_, 
        stg2_real_2__0_}) );
  FFT_ultrafast2_shift_DW01_add_10 add_311 ( .A({stg1_real_1__15_, 
        stg1_real_1__14_, stg1_real_1__13_, stg1_real_1__12_, stg1_real_1__11_, 
        stg1_real_1__10_, stg1_real_1__9_, stg1_real_1__8_, stg1_real_1__7_, 
        stg1_real_1__6_, stg1_real_1__5_, stg1_real_1__4_, stg1_real_1__3_, 
        stg1_real_1__2_, stg1_real_1__1_, stg1_real_1__0_}), .B({
        stg1_real_5__15_, stg1_real_5__14_, stg1_real_5__13_, stg1_real_5__12_, 
        stg1_real_5__11_, stg1_real_5__10_, stg1_real_5__9_, stg1_real_5__8_, 
        stg1_real_5__7_, stg1_real_5__6_, stg1_real_5__5_, stg1_real_5__4_, 
        stg1_real_5__3_, stg1_real_5__2_, stg1_real_5__1_, stg1_real_5__0_}), 
        .SUM({stg2_real_1__15_, stg2_real_1__14_, stg2_real_1__13_, 
        stg2_real_1__12_, stg2_real_1__11_, stg2_real_1__10_, stg2_real_1__9_, 
        stg2_real_1__8_, stg2_real_1__7_, stg2_real_1__6_, stg2_real_1__5_, 
        stg2_real_1__4_, stg2_real_1__3_, stg2_real_1__2_, stg2_real_1__1_, 
        stg2_real_1__0_}) );
  FFT_ultrafast2_shift_DW01_add_11 add_310 ( .A({stg1_real_0__15_, 
        stg1_real_0__14_, stg1_real_0__13_, stg1_real_0__12_, stg1_real_0__11_, 
        stg1_real_0__10_, stg1_real_0__9_, stg1_real_0__8_, stg1_real_0__7_, 
        stg1_real_0__6_, stg1_real_0__5_, stg1_real_0__4_, stg1_real_0__3_, 
        stg1_real_0__2_, stg1_real_0__1_, stg1_real_0__0_}), .B({
        stg1_real_4__15_, stg1_real_4__14_, stg1_real_4__13_, stg1_real_4__12_, 
        stg1_real_4__11_, stg1_real_4__10_, stg1_real_4__9_, stg1_real_4__8_, 
        stg1_real_4__7_, stg1_real_4__6_, stg1_real_4__5_, stg1_real_4__4_, 
        stg1_real_4__3_, stg1_real_4__2_, stg1_real_4__1_, stg1_real_4__0_}), 
        .SUM({stg2_real_0__15_, stg2_real_0__14_, stg2_real_0__13_, 
        stg2_real_0__12_, stg2_real_0__11_, stg2_real_0__10_, stg2_real_0__9_, 
        stg2_real_0__8_, stg2_real_0__7_, stg2_real_0__6_, stg2_real_0__5_, 
        stg2_real_0__4_, stg2_real_0__3_, stg2_real_0__2_, stg2_real_0__1_, 
        stg2_real_0__0_}) );
  FFT_ultrafast2_shift_DW01_sub_16 sub_308 ( .A(fir_d), .B({data_7__15_, 
        data_7__14_, data_7__13_, data_7__12_, data_7__11_, data_7__10_, 
        data_7__9_, data_7__8_, data_7__7_, data_7__6_, data_7__5_, data_7__4_, 
        data_7__3_, data_7__2_, data_7__1_, data_7__0_}), .DIFF({
        stg2_img_11__15_, stg2_img_11__14_, stg2_img_11__13_, stg2_img_11__12_, 
        stg2_img_11__11_, stg2_img_11__10_, stg2_img_11__9_, stg2_img_11__8_, 
        stg2_img_11__7_, stg2_img_11__6_, stg2_img_11__5_, stg2_img_11__4_, 
        stg2_img_11__3_, stg2_img_11__2_, stg2_img_11__1_, stg2_img_15__0_})
         );
  FFT_ultrafast2_shift_DW01_sub_17 sub_307 ( .A({data_14__15_, data_14__14_, 
        data_14__13_, data_14__12_, data_14__11_, data_14__10_, data_14__9_, 
        data_14__8_, data_14__7_, data_14__6_, data_14__5_, data_14__4_, 
        data_14__3_, data_14__2_, data_14__1_, data_14__0_}), .B({data_6__15_, 
        data_6__14_, data_6__13_, data_6__12_, data_6__11_, data_6__10_, 
        data_6__9_, data_6__8_, data_6__7_, data_6__6_, data_6__5_, data_6__4_, 
        data_6__3_, data_6__2_, data_6__1_, data_6__0_}), .DIFF({
        stg2_img_10__15_, stg2_img_10__14_, stg2_img_10__13_, stg2_img_10__12_, 
        stg2_img_10__11_, stg2_img_10__10_, stg2_img_10__9_, stg2_img_10__8_, 
        stg2_img_10__7_, stg2_img_10__6_, stg2_img_10__5_, stg2_img_10__4_, 
        stg2_img_10__3_, stg2_img_10__2_, stg2_img_10__1_, stg2_img_14__0_})
         );
  FFT_ultrafast2_shift_DW01_sub_18 sub_306 ( .A({data_13__15_, data_13__14_, 
        data_13__13_, data_13__12_, data_13__11_, data_13__10_, data_13__9_, 
        data_13__8_, data_13__7_, data_13__6_, data_13__5_, data_13__4_, 
        data_13__3_, data_13__2_, data_13__1_, data_13__0_}), .B({data_5__15_, 
        data_5__14_, data_5__13_, data_5__12_, data_5__11_, data_5__10_, 
        data_5__9_, data_5__8_, data_5__7_, data_5__6_, data_5__5_, data_5__4_, 
        data_5__3_, data_5__2_, data_5__1_, data_5__0_}), .DIFF({
        stg2_img_9__15_, stg2_img_9__14_, stg2_img_9__13_, stg2_img_9__12_, 
        stg2_img_9__11_, stg2_img_9__10_, stg2_img_9__9_, stg2_img_9__8_, 
        stg2_img_9__7_, stg2_img_9__6_, stg2_img_9__5_, stg2_img_9__4_, 
        stg2_img_9__3_, stg2_img_9__2_, stg2_img_9__1_, stg2_img_13__0_}) );
  FFT_ultrafast2_shift_DW01_sub_19 sub_305 ( .A({data_12__15_, data_12__14_, 
        data_12__13_, data_12__12_, data_12__11_, data_12__10_, data_12__9_, 
        data_12__8_, data_12__7_, data_12__6_, data_12__5_, data_12__4_, 
        data_12__3_, data_12__2_, data_12__1_, data_12__0_}), .B({data_4__15_, 
        data_4__14_, data_4__13_, data_4__12_, data_4__11_, data_4__10_, 
        data_4__9_, data_4__8_, data_4__7_, data_4__6_, data_4__5_, data_4__4_, 
        data_4__3_, data_4__2_, data_4__1_, data_4__0_}), .DIFF({
        stg2_img_8__15_, stg2_img_8__14_, stg2_img_8__13_, stg2_img_8__12_, 
        stg2_img_8__11_, stg2_img_8__10_, stg2_img_8__9_, stg2_img_8__8_, 
        stg2_img_8__7_, stg2_img_8__6_, stg2_img_8__5_, stg2_img_8__4_, 
        stg2_img_8__3_, stg2_img_8__2_, stg2_img_8__1_, stg2_img_8__0_}) );
  FFT_ultrafast2_shift_DW01_sub_20 sub_287 ( .A({data_3__15_, data_3__14_, 
        data_3__13_, data_3__12_, data_3__11_, data_3__10_, data_3__9_, 
        data_3__8_, data_3__7_, data_3__6_, data_3__5_, data_3__4_, data_3__3_, 
        data_3__2_, data_3__1_, data_3__0_}), .B({data_11__15_, data_11__14_, 
        data_11__13_, data_11__12_, data_11__11_, data_11__10_, data_11__9_, 
        data_11__8_, data_11__7_, data_11__6_, data_11__5_, data_11__4_, 
        data_11__3_, data_11__2_, data_11__1_, data_11__0_}), .DIFF({
        stg2_real_15__15_, stg2_real_15__14_, stg2_real_15__13_, 
        stg2_real_15__12_, stg2_real_15__11_, stg2_real_15__10_, 
        stg2_real_15__9_, stg2_real_15__8_, stg2_real_15__7_, stg2_real_15__6_, 
        stg2_real_15__5_, stg2_real_15__4_, stg2_real_15__3_, stg2_real_15__2_, 
        stg2_real_15__1_, stg2_real_15__0_}) );
  FFT_ultrafast2_shift_DW01_sub_21 sub_286 ( .A({data_2__15_, data_2__14_, 
        data_2__13_, data_2__12_, data_2__11_, data_2__10_, data_2__9_, 
        data_2__8_, data_2__7_, data_2__6_, data_2__5_, data_2__4_, data_2__3_, 
        data_2__2_, data_2__1_, data_2__0_}), .B({data_10__15_, data_10__14_, 
        data_10__13_, data_10__12_, data_10__11_, data_10__10_, data_10__9_, 
        data_10__8_, data_10__7_, data_10__6_, data_10__5_, data_10__4_, 
        data_10__3_, data_10__2_, data_10__1_, data_10__0_}), .DIFF({
        stg2_real_14__15_, stg2_real_14__14_, stg2_real_14__13_, 
        stg2_real_14__12_, stg2_real_14__11_, stg2_real_14__10_, 
        stg2_real_14__9_, stg2_real_14__8_, stg2_real_14__7_, stg2_real_14__6_, 
        stg2_real_14__5_, stg2_real_14__4_, stg2_real_14__3_, stg2_real_14__2_, 
        stg2_real_14__1_, stg2_real_14__0_}) );
  FFT_ultrafast2_shift_DW01_sub_22 sub_285 ( .A({data_1__15_, data_1__14_, 
        data_1__13_, data_1__12_, data_1__11_, data_1__10_, data_1__9_, 
        data_1__8_, data_1__7_, data_1__6_, data_1__5_, data_1__4_, data_1__3_, 
        data_1__2_, data_1__1_, data_1__0_}), .B({data_9__15_, data_9__14_, 
        data_9__13_, data_9__12_, data_9__11_, data_9__10_, data_9__9_, 
        data_9__8_, data_9__7_, data_9__6_, data_9__5_, data_9__4_, data_9__3_, 
        data_9__2_, data_9__1_, data_9__0_}), .DIFF({stg2_real_13__15_, 
        stg2_real_13__14_, stg2_real_13__13_, stg2_real_13__12_, 
        stg2_real_13__11_, stg2_real_13__10_, stg2_real_13__9_, 
        stg2_real_13__8_, stg2_real_13__7_, stg2_real_13__6_, stg2_real_13__5_, 
        stg2_real_13__4_, stg2_real_13__3_, stg2_real_13__2_, stg2_real_13__1_, 
        stg2_real_13__0_}) );
  FFT_ultrafast2_shift_DW01_sub_23 sub_284 ( .A({data_0__15_, data_0__14_, 
        data_0__13_, data_0__12_, data_0__11_, data_0__10_, data_0__9_, 
        data_0__8_, data_0__7_, data_0__6_, data_0__5_, data_0__4_, data_0__3_, 
        data_0__2_, data_0__1_, data_0__0_}), .B({data_8__15_, data_8__14_, 
        data_8__13_, data_8__12_, data_8__11_, data_8__10_, data_8__9_, 
        data_8__8_, data_8__7_, data_8__6_, data_8__5_, data_8__4_, data_8__3_, 
        data_8__2_, data_8__1_, data_8__0_}), .DIFF({stg2_real_12__15_, 
        stg2_real_12__14_, stg2_real_12__13_, stg2_real_12__12_, 
        stg2_real_12__11_, stg2_real_12__10_, stg2_real_12__9_, 
        stg2_real_12__8_, stg2_real_12__7_, stg2_real_12__6_, stg2_real_12__5_, 
        stg2_real_12__4_, stg2_real_12__3_, stg2_real_12__2_, stg2_real_12__1_, 
        stg2_real_12__0_}) );
  FFT_ultrafast2_shift_DW01_add_12 add_283 ( .A({data_7__15_, data_7__14_, 
        data_7__13_, data_7__12_, data_7__11_, data_7__10_, data_7__9_, 
        data_7__8_, data_7__7_, data_7__6_, data_7__5_, data_7__4_, data_7__3_, 
        data_7__2_, data_7__1_, data_7__0_}), .B(fir_d), .SUM({
        stg1_real_7__15_, stg1_real_7__14_, stg1_real_7__13_, stg1_real_7__12_, 
        stg1_real_7__11_, stg1_real_7__10_, stg1_real_7__9_, stg1_real_7__8_, 
        stg1_real_7__7_, stg1_real_7__6_, stg1_real_7__5_, stg1_real_7__4_, 
        stg1_real_7__3_, stg1_real_7__2_, stg1_real_7__1_, stg1_real_7__0_})
         );
  FFT_ultrafast2_shift_DW01_add_13 add_282 ( .A({data_6__15_, data_6__14_, 
        data_6__13_, data_6__12_, data_6__11_, data_6__10_, data_6__9_, 
        data_6__8_, data_6__7_, data_6__6_, data_6__5_, data_6__4_, data_6__3_, 
        data_6__2_, data_6__1_, data_6__0_}), .B({data_14__15_, data_14__14_, 
        data_14__13_, data_14__12_, data_14__11_, data_14__10_, data_14__9_, 
        data_14__8_, data_14__7_, data_14__6_, data_14__5_, data_14__4_, 
        data_14__3_, data_14__2_, data_14__1_, data_14__0_}), .SUM({
        stg1_real_6__15_, stg1_real_6__14_, stg1_real_6__13_, stg1_real_6__12_, 
        stg1_real_6__11_, stg1_real_6__10_, stg1_real_6__9_, stg1_real_6__8_, 
        stg1_real_6__7_, stg1_real_6__6_, stg1_real_6__5_, stg1_real_6__4_, 
        stg1_real_6__3_, stg1_real_6__2_, stg1_real_6__1_, stg1_real_6__0_})
         );
  FFT_ultrafast2_shift_DW01_add_14 add_281 ( .A({data_5__15_, data_5__14_, 
        data_5__13_, data_5__12_, data_5__11_, data_5__10_, data_5__9_, 
        data_5__8_, data_5__7_, data_5__6_, data_5__5_, data_5__4_, data_5__3_, 
        data_5__2_, data_5__1_, data_5__0_}), .B({data_13__15_, data_13__14_, 
        data_13__13_, data_13__12_, data_13__11_, data_13__10_, data_13__9_, 
        data_13__8_, data_13__7_, data_13__6_, data_13__5_, data_13__4_, 
        data_13__3_, data_13__2_, data_13__1_, data_13__0_}), .SUM({
        stg1_real_5__15_, stg1_real_5__14_, stg1_real_5__13_, stg1_real_5__12_, 
        stg1_real_5__11_, stg1_real_5__10_, stg1_real_5__9_, stg1_real_5__8_, 
        stg1_real_5__7_, stg1_real_5__6_, stg1_real_5__5_, stg1_real_5__4_, 
        stg1_real_5__3_, stg1_real_5__2_, stg1_real_5__1_, stg1_real_5__0_})
         );
  FFT_ultrafast2_shift_DW01_add_15 add_280 ( .A({data_4__15_, data_4__14_, 
        data_4__13_, data_4__12_, data_4__11_, data_4__10_, data_4__9_, 
        data_4__8_, data_4__7_, data_4__6_, data_4__5_, data_4__4_, data_4__3_, 
        data_4__2_, data_4__1_, data_4__0_}), .B({data_12__15_, data_12__14_, 
        data_12__13_, data_12__12_, data_12__11_, data_12__10_, data_12__9_, 
        data_12__8_, data_12__7_, data_12__6_, data_12__5_, data_12__4_, 
        data_12__3_, data_12__2_, data_12__1_, data_12__0_}), .SUM({
        stg1_real_4__15_, stg1_real_4__14_, stg1_real_4__13_, stg1_real_4__12_, 
        stg1_real_4__11_, stg1_real_4__10_, stg1_real_4__9_, stg1_real_4__8_, 
        stg1_real_4__7_, stg1_real_4__6_, stg1_real_4__5_, stg1_real_4__4_, 
        stg1_real_4__3_, stg1_real_4__2_, stg1_real_4__1_, stg1_real_4__0_})
         );
  FFT_ultrafast2_shift_DW01_add_16 add_279 ( .A({data_3__15_, data_3__14_, 
        data_3__13_, data_3__12_, data_3__11_, data_3__10_, data_3__9_, 
        data_3__8_, data_3__7_, data_3__6_, data_3__5_, data_3__4_, data_3__3_, 
        data_3__2_, data_3__1_, data_3__0_}), .B({data_11__15_, data_11__14_, 
        data_11__13_, data_11__12_, data_11__11_, data_11__10_, data_11__9_, 
        data_11__8_, data_11__7_, data_11__6_, data_11__5_, data_11__4_, 
        data_11__3_, data_11__2_, data_11__1_, data_11__0_}), .SUM({
        stg1_real_3__15_, stg1_real_3__14_, stg1_real_3__13_, stg1_real_3__12_, 
        stg1_real_3__11_, stg1_real_3__10_, stg1_real_3__9_, stg1_real_3__8_, 
        stg1_real_3__7_, stg1_real_3__6_, stg1_real_3__5_, stg1_real_3__4_, 
        stg1_real_3__3_, stg1_real_3__2_, stg1_real_3__1_, stg1_real_3__0_})
         );
  FFT_ultrafast2_shift_DW01_add_17 add_278 ( .A({data_2__15_, data_2__14_, 
        data_2__13_, data_2__12_, data_2__11_, data_2__10_, data_2__9_, 
        data_2__8_, data_2__7_, data_2__6_, data_2__5_, data_2__4_, data_2__3_, 
        data_2__2_, data_2__1_, data_2__0_}), .B({data_10__15_, data_10__14_, 
        data_10__13_, data_10__12_, data_10__11_, data_10__10_, data_10__9_, 
        data_10__8_, data_10__7_, data_10__6_, data_10__5_, data_10__4_, 
        data_10__3_, data_10__2_, data_10__1_, data_10__0_}), .SUM({
        stg1_real_2__15_, stg1_real_2__14_, stg1_real_2__13_, stg1_real_2__12_, 
        stg1_real_2__11_, stg1_real_2__10_, stg1_real_2__9_, stg1_real_2__8_, 
        stg1_real_2__7_, stg1_real_2__6_, stg1_real_2__5_, stg1_real_2__4_, 
        stg1_real_2__3_, stg1_real_2__2_, stg1_real_2__1_, stg1_real_2__0_})
         );
  FFT_ultrafast2_shift_DW01_add_18 add_277 ( .A({data_1__15_, data_1__14_, 
        data_1__13_, data_1__12_, data_1__11_, data_1__10_, data_1__9_, 
        data_1__8_, data_1__7_, data_1__6_, data_1__5_, data_1__4_, data_1__3_, 
        data_1__2_, data_1__1_, data_1__0_}), .B({data_9__15_, data_9__14_, 
        data_9__13_, data_9__12_, data_9__11_, data_9__10_, data_9__9_, 
        data_9__8_, data_9__7_, data_9__6_, data_9__5_, data_9__4_, data_9__3_, 
        data_9__2_, data_9__1_, data_9__0_}), .SUM({stg1_real_1__15_, 
        stg1_real_1__14_, stg1_real_1__13_, stg1_real_1__12_, stg1_real_1__11_, 
        stg1_real_1__10_, stg1_real_1__9_, stg1_real_1__8_, stg1_real_1__7_, 
        stg1_real_1__6_, stg1_real_1__5_, stg1_real_1__4_, stg1_real_1__3_, 
        stg1_real_1__2_, stg1_real_1__1_, stg1_real_1__0_}) );
  FFT_ultrafast2_shift_DW01_add_19 add_276 ( .A({data_0__15_, data_0__14_, 
        data_0__13_, data_0__12_, data_0__11_, data_0__10_, data_0__9_, 
        data_0__8_, data_0__7_, data_0__6_, data_0__5_, data_0__4_, data_0__3_, 
        data_0__2_, data_0__1_, data_0__0_}), .B({data_8__15_, data_8__14_, 
        data_8__13_, data_8__12_, data_8__11_, data_8__10_, data_8__9_, 
        data_8__8_, data_8__7_, data_8__6_, data_8__5_, data_8__4_, data_8__3_, 
        data_8__2_, data_8__1_, data_8__0_}), .SUM({stg1_real_0__15_, 
        stg1_real_0__14_, stg1_real_0__13_, stg1_real_0__12_, stg1_real_0__11_, 
        stg1_real_0__10_, stg1_real_0__9_, stg1_real_0__8_, stg1_real_0__7_, 
        stg1_real_0__6_, stg1_real_0__5_, stg1_real_0__4_, stg1_real_0__3_, 
        stg1_real_0__2_, stg1_real_0__1_, stg1_real_0__0_}) );
  FFT_ultrafast2_shift_DW_mult_uns_8 mult_232 ( .a_15_(mul_2_in[15]), .a_14_(
        mul_2_in[14]), .a_13_(mul_2_in[13]), .a_12_(mul_2_in[12]), .a_11_(
        mul_2_in[11]), .a_10_(mul_2_in[10]), .a_9_(mul_2_in[9]), .a_8_(
        mul_2_in[8]), .a_7_(mul_2_in[7]), .a_6_(mul_2_in[6]), .a_5_(
        mul_2_in[5]), .a_4_(mul_2_in[4]), .a_3_(mul_2_in[3]), .a_2_(
        mul_2_in[2]), .a_1_(n212), .a_0_(mul_2_in[0]), .b_31_(mul_0_Wn_19), 
        .b_30_(mul_0_Wn_19), .b_29_(mul_0_Wn_19), .b_28_(mul_0_Wn_19), .b_27_(
        mul_0_Wn_19), .b_26_(mul_0_Wn_19), .b_25_(mul_0_Wn_19), .b_16_(
        mul_0_Wn_19), .b_15_(mul_0_Wn[15]), .b_14_(n88), .b_13_(mul_0_Wn[13]), 
        .b_12_(mul_0_Wn[12]), .b_11_(mul_0_Wn[11]), .b_10_(mul_0_Wn[15]), 
        .b_9_(mul_0_Wn_19), .b_8_(mul_0_Wn_8), .b_7_(n88), .b_6_(mul_0_Wn_6), 
        .b_5_(mul_0_Wn_6), .b_4_(mul_0_Wn_6), .b_3_(mul_0_Wn_19), .b_2_(n86), 
        .b_1_(n85), .b_0_(mul_0_Wn_0), .product_31_(mul_0_out_31_), 
        .product_30_(mul_0_out_30_), .product_29_(mul_0_out_29_), 
        .product_28_(mul_0_out_28_), .product_27_(mul_0_out_27_), 
        .product_26_(mul_0_out_26_), .product_25_(mul_0_out_25_), 
        .product_24_(mul_0_out_24_), .product_23_(mul_0_out_23_), 
        .product_22_(mul_0_out_22_), .product_21_(mul_0_out_21_), 
        .product_20_(mul_0_out_20_), .product_19_(mul_0_out_19_), 
        .product_18_(mul_0_out_18_), .product_17_(mul_0_out_17_), 
        .product_16_(mul_0_out_16_), .product_15_(mul_0_out_15_), 
        .product_14_(mul_0_out_14_), .product_13_(mul_0_out_13_), 
        .product_12_(mul_0_out_12_), .product_11_(mul_0_out_11_), 
        .product_10_(mul_0_out_10_), .product_9_(mul_0_out_9_), .product_8_(
        mul_0_out_8_), .product_7_(mul_0_out_7_), .product_6_(mul_0_out_6_), 
        .product_5_(mul_0_out_5_), .product_4_(mul_0_out_4_), .product_3_(
        mul_0_out_3_), .product_2_(mul_0_out_2_), .product_1_(mul_0_out_1_), 
        .product_0_(mul_0_out_0_) );
  FFT_ultrafast2_shift_DW_mult_uns_9 mult_250 ( .a_15_(mul_1_in[15]), .a_14_(
        mul_1_in[14]), .a_13_(mul_1_in[13]), .a_12_(mul_1_in[12]), .a_11_(
        mul_1_in[11]), .a_10_(mul_1_in[10]), .a_9_(mul_1_in[9]), .a_8_(
        mul_1_in[8]), .a_7_(mul_1_in[7]), .a_6_(mul_1_in[6]), .a_5_(
        mul_1_in[5]), .a_4_(mul_1_in[4]), .a_3_(mul_1_in[3]), .a_2_(
        mul_1_in[2]), .a_1_(mul_1_in[1]), .a_0_(mul_1_in[0]), .b_16_(
        mul_0_Wn_19), .b_15_(mul_0_Wn[15]), .b_14_(n88), .b_13_(mul_0_Wn[13]), 
        .b_12_(mul_0_Wn[12]), .b_11_(mul_0_Wn[11]), .b_10_(mul_0_Wn[15]), 
        .b_9_(mul_0_Wn_19), .b_8_(mul_0_Wn_8), .b_7_(n88), .b_6_(mul_0_Wn_6), 
        .b_5_(mul_0_Wn_6), .b_4_(mul_0_Wn_6), .b_3_(mul_0_Wn_19), .b_2_(n87), 
        .b_1_(n85), .b_0_(mul_0_Wn_0), .product_31_(mul_3_out_31_), 
        .product_30_(mul_3_out_30_), .product_29_(mul_3_out_29_), 
        .product_28_(mul_3_out_28_), .product_27_(mul_3_out_27_), 
        .product_26_(mul_3_out_26_), .product_25_(mul_3_out_25_), 
        .product_24_(mul_3_out_24_), .product_23_(mul_3_out_23_), 
        .product_22_(mul_3_out_22_), .product_21_(mul_3_out_21_), 
        .product_20_(mul_3_out_20_), .product_19_(mul_3_out_19_), 
        .product_18_(mul_3_out_18_), .product_17_(mul_3_out_17_), 
        .product_16_(mul_3_out_16_), .product_15_(mul_3_out_15_), 
        .product_14_(mul_3_out_14_), .product_13_(mul_3_out_13_), 
        .product_12_(mul_3_out_12_), .product_11_(mul_3_out_11_), 
        .product_10_(mul_3_out_10_), .product_9_(mul_3_out_9_), .product_8_(
        mul_3_out_8_), .product_7_(mul_3_out_7_), .product_6_(mul_3_out_6_), 
        .product_5_(mul_3_out_5_), .product_4_(mul_3_out_4_), .product_3_(
        mul_3_out_3_), .product_2_(mul_3_out_2_), .product_1_(mul_3_out_1_), 
        .product_0_(mul_3_out_0_) );
  FFT_ultrafast2_shift_DW_mult_uns_10 mult_245 ( .a_15_(mul_2_in[15]), .a_14_(
        mul_2_in[14]), .a_13_(mul_2_in[13]), .a_12_(mul_2_in[12]), .a_11_(
        mul_2_in[11]), .a_10_(mul_2_in[10]), .a_9_(mul_2_in[9]), .a_8_(
        mul_2_in[8]), .a_7_(mul_2_in[7]), .a_6_(mul_2_in[6]), .a_5_(
        mul_2_in[5]), .a_4_(mul_2_in[4]), .a_3_(mul_2_in[3]), .a_2_(
        mul_2_in[2]), .a_1_(n212), .a_0_(mul_2_in[0]), .b_16_(mul_2_Wn_19), 
        .b_15_(n209), .b_14_(mul_2_Wn[14]), .b_13_(mul_2_Wn[13]), .b_12_(n85), 
        .b_11_(mul_2_Wn_11), .b_10_(n209), .b_9_(mul_2_Wn_9), .b_8_(mul_2_Wn_8), .b_7_(mul_2_Wn[14]), .b_6_(n87), .b_5_(n87), .b_4_(n87), .b_3_(mul_2_Wn_9), 
        .b_2_(n86), .b_1_(n10370), .b_0_(mul_0_Wn_0), .product_31_(
        mul_2_out_31_), .product_30_(mul_2_out_30_), .product_29_(
        mul_2_out_29_), .product_28_(mul_2_out_28_), .product_27_(
        mul_2_out_27_), .product_26_(mul_2_out_26_), .product_25_(
        mul_2_out_25_), .product_24_(mul_2_out_24_), .product_23_(
        mul_2_out_23_), .product_22_(mul_2_out_22_), .product_21_(
        mul_2_out_21_), .product_20_(mul_2_out_20_), .product_19_(
        mul_2_out_19_), .product_18_(mul_2_out_18_), .product_17_(
        mul_2_out_17_), .product_16_(mul_2_out_16_), .product_15_(
        mul_2_out_15_), .product_14_(mul_2_out_14_), .product_13_(
        mul_2_out_13_), .product_12_(mul_2_out_12_), .product_11_(
        mul_2_out_11_), .product_10_(mul_2_out_10_), .product_9_(mul_2_out_9_), 
        .product_8_(mul_2_out_8_), .product_7_(mul_2_out_7_), .product_6_(
        mul_2_out_6_), .product_5_(mul_2_out_5_), .product_4_(mul_2_out_4_), 
        .product_3_(mul_2_out_3_), .product_2_(mul_2_out_2_), .product_1_(
        mul_2_out_1_), .product_0_(mul_2_out_0_) );
  FFT_ultrafast2_shift_DW01_add_22 add_253 ( .A({mul_2_out_31_, mul_2_out_30_, 
        mul_2_out_29_, mul_2_out_28_, mul_2_out_27_, mul_2_out_26_, 
        mul_2_out_25_, mul_2_out_24_, mul_2_out_23_, mul_2_out_22_, 
        mul_2_out_21_, mul_2_out_20_, mul_2_out_19_, mul_2_out_18_, 
        mul_2_out_17_, mul_2_out_16_, mul_2_out_15_, mul_2_out_14_, 
        mul_2_out_13_, mul_2_out_12_, mul_2_out_11_, mul_2_out_10_, 
        mul_2_out_9_, mul_2_out_8_, mul_2_out_7_, mul_2_out_6_, mul_2_out_5_, 
        mul_2_out_4_, mul_2_out_3_, mul_2_out_2_, mul_2_out_1_, mul_2_out_0_}), 
        .B({mul_3_out_31_, mul_3_out_30_, mul_3_out_29_, mul_3_out_28_, 
        mul_3_out_27_, mul_3_out_26_, mul_3_out_25_, mul_3_out_24_, 
        mul_3_out_23_, mul_3_out_22_, mul_3_out_21_, mul_3_out_20_, 
        mul_3_out_19_, mul_3_out_18_, mul_3_out_17_, mul_3_out_16_, 
        mul_3_out_15_, mul_3_out_14_, mul_3_out_13_, mul_3_out_12_, 
        mul_3_out_11_, mul_3_out_10_, mul_3_out_9_, mul_3_out_8_, mul_3_out_7_, 
        mul_3_out_6_, mul_3_out_5_, mul_3_out_4_, mul_3_out_3_, mul_3_out_2_, 
        mul_3_out_1_, mul_3_out_0_}), .SUM_31_(mul_o_add[31]), .SUM_30_(
        mul_o_add[30]), .SUM_29_(mul_o_add[29]), .SUM_28_(mul_o_add[28]), 
        .SUM_27_(mul_o_add[27]), .SUM_26_(mul_o_add[26]), .SUM_25_(
        mul_o_add[25]), .SUM_24_(mul_o_add[24]), .SUM_23_(mul_o_add[23]), 
        .SUM_22_(mul_o_add[22]), .SUM_21_(mul_o_add[21]), .SUM_20_(
        mul_o_add[20]), .SUM_19_(mul_o_add[19]), .SUM_18_(mul_o_add[18]), 
        .SUM_17_(mul_o_add[17]), .SUM_16_(mul_o_add[16]) );
  FFT_ultrafast2_shift_DW_mult_uns_11 mult_237 ( .a_15_(mul_1_in[15]), .a_14_(
        mul_1_in[14]), .a_13_(mul_1_in[13]), .a_12_(mul_1_in[12]), .a_11_(
        mul_1_in[11]), .a_10_(mul_1_in[10]), .a_9_(mul_1_in[9]), .a_8_(
        mul_1_in[8]), .a_7_(mul_1_in[7]), .a_6_(mul_1_in[6]), .a_5_(
        mul_1_in[5]), .a_4_(mul_1_in[4]), .a_3_(mul_1_in[3]), .a_2_(
        mul_1_in[2]), .a_1_(mul_1_in[1]), .a_0_(mul_1_in[0]), .b_16_(
        mul_2_Wn_19), .b_15_(n209), .b_14_(mul_2_Wn[14]), .b_13_(mul_2_Wn[13]), 
        .b_12_(n85), .b_11_(mul_2_Wn_11), .b_10_(n209), .b_9_(mul_2_Wn_9), 
        .b_8_(mul_2_Wn_8), .b_7_(mul_2_Wn[14]), .b_6_(n87), .b_5_(n87), .b_4_(
        n87), .b_3_(mul_2_Wn_9), .b_2_(n87), .b_1_(mul_2_Wn[13]), .b_0_(
        mul_0_Wn_0), .product_31_(mul_1_out_31_), .product_30_(mul_1_out_30_), 
        .product_29_(mul_1_out_29_), .product_28_(mul_1_out_28_), 
        .product_27_(mul_1_out_27_), .product_26_(mul_1_out_26_), 
        .product_25_(mul_1_out_25_), .product_24_(mul_1_out_24_), 
        .product_23_(mul_1_out_23_), .product_22_(mul_1_out_22_), 
        .product_21_(mul_1_out_21_), .product_20_(mul_1_out_20_), 
        .product_19_(mul_1_out_19_), .product_18_(mul_1_out_18_), 
        .product_17_(mul_1_out_17_), .product_16_(mul_1_out_16_), 
        .product_15_(mul_1_out_15_), .product_14_(mul_1_out_14_), 
        .product_13_(mul_1_out_13_), .product_12_(mul_1_out_12_), 
        .product_11_(mul_1_out_11_), .product_10_(mul_1_out_10_), .product_9_(
        mul_1_out_9_), .product_8_(mul_1_out_8_), .product_7_(mul_1_out_7_), 
        .product_6_(mul_1_out_6_), .product_5_(mul_1_out_5_), .product_4_(
        mul_1_out_4_), .product_3_(mul_1_out_3_), .product_2_(mul_1_out_2_), 
        .product_1_(mul_1_out_1_), .product_0_(mul_1_out_0_) );
  FFT_ultrafast2_shift_DW01_sub_26 sub_240 ( .A({mul_0_out_31_, mul_0_out_30_, 
        mul_0_out_29_, mul_0_out_28_, mul_0_out_27_, mul_0_out_26_, 
        mul_0_out_25_, mul_0_out_24_, mul_0_out_23_, mul_0_out_22_, 
        mul_0_out_21_, mul_0_out_20_, mul_0_out_19_, mul_0_out_18_, 
        mul_0_out_17_, mul_0_out_16_, mul_0_out_15_, mul_0_out_14_, 
        mul_0_out_13_, mul_0_out_12_, mul_0_out_11_, mul_0_out_10_, 
        mul_0_out_9_, mul_0_out_8_, mul_0_out_7_, mul_0_out_6_, mul_0_out_5_, 
        mul_0_out_4_, mul_0_out_3_, mul_0_out_2_, mul_0_out_1_, mul_0_out_0_}), 
        .B({mul_1_out_31_, mul_1_out_30_, mul_1_out_29_, mul_1_out_28_, 
        mul_1_out_27_, mul_1_out_26_, mul_1_out_25_, mul_1_out_24_, 
        mul_1_out_23_, mul_1_out_22_, mul_1_out_21_, mul_1_out_20_, 
        mul_1_out_19_, mul_1_out_18_, mul_1_out_17_, mul_1_out_16_, 
        mul_1_out_15_, mul_1_out_14_, mul_1_out_13_, mul_1_out_12_, 
        mul_1_out_11_, mul_1_out_10_, mul_1_out_9_, mul_1_out_8_, mul_1_out_7_, 
        mul_1_out_6_, mul_1_out_5_, mul_1_out_4_, mul_1_out_3_, mul_1_out_2_, 
        mul_1_out_1_, mul_1_out_0_}), .DIFF_31_(mul_o_sub[31]), .DIFF_30_(
        mul_o_sub[30]), .DIFF_29_(mul_o_sub[29]), .DIFF_28_(mul_o_sub[28]), 
        .DIFF_27_(mul_o_sub[27]), .DIFF_26_(mul_o_sub[26]), .DIFF_25_(
        mul_o_sub[25]), .DIFF_24_(mul_o_sub[24]), .DIFF_23_(mul_o_sub[23]), 
        .DIFF_22_(mul_o_sub[22]), .DIFF_21_(mul_o_sub[21]), .DIFF_20_(
        mul_o_sub[20]), .DIFF_19_(mul_o_sub[19]), .DIFF_18_(mul_o_sub[18]), 
        .DIFF_17_(mul_o_sub[17]), .DIFF_16_(mul_o_sub[16]) );
  DFFRX1 first_cnt_reg ( .D(n1792), .CK(clk), .RN(n3149), .QN(n1791) );
  DFFQX1 data_reg_0__15_ ( .D(data_1__15_), .CK(clk), .Q(data_0__15_) );
  DFFQX1 data_reg_8__15_ ( .D(data_9__15_), .CK(clk), .Q(data_8__15_) );
  DFFQX1 stg_reg_reg_4__28_ ( .D(n3212), .CK(clk), .Q(stg_reg[156]) );
  DFFQX1 stg_reg_reg_4__29_ ( .D(n3211), .CK(clk), .Q(stg_reg[157]) );
  DFFQX1 stg_reg_reg_4__30_ ( .D(n3210), .CK(clk), .Q(stg_reg[158]) );
  DFFQX1 stg_reg_reg_4__31_ ( .D(n3209), .CK(clk), .Q(stg_reg[159]) );
  DFFX1 stg_reg_reg_3__30_ ( .D(n2277), .CK(clk), .Q(n1767), .QN(n2567) );
  DFFX1 stg_reg_reg_3__31_ ( .D(n2276), .CK(clk), .Q(n1769), .QN(n2559) );
  DFFX1 stg_reg_reg_12__28_ ( .D(n2119), .CK(clk), .Q(n1624), .QN(n1175) );
  DFFX1 stg_reg_reg_12__29_ ( .D(n2118), .CK(clk), .Q(n1627), .QN(n1166) );
  DFFX1 stg_reg_reg_8__29_ ( .D(n2150), .CK(clk), .Q(n1626), .QN(n1165) );
  DFFX1 stg_reg_reg_0__29_ ( .D(n2182), .CK(clk), .Q(n1625), .QN(n1162) );
  DFFX1 stg_reg_reg_12__30_ ( .D(n2117), .CK(clk), .Q(n1630), .QN(n1157) );
  DFFX1 stg_reg_reg_8__30_ ( .D(n2149), .CK(clk), .Q(n1629), .QN(n1156) );
  DFFX1 stg_reg_reg_0__30_ ( .D(n2181), .CK(clk), .Q(n1628), .QN(n1153) );
  DFFX1 stg_reg_reg_12__31_ ( .D(n2116), .CK(clk), .Q(n1633), .QN(n2707) );
  DFFX1 stg_reg_reg_8__31_ ( .D(n2148), .CK(clk), .Q(n1632), .QN(n2706) );
  DFFX1 stg_reg_reg_0__31_ ( .D(n2180), .CK(clk), .Q(n1631), .QN(n2703) );
  DFFX1 stg_reg_reg_2__30_ ( .D(n2245), .CK(clk), .Q(n1724), .QN(n1295) );
  DFFX1 stg_reg_reg_2__31_ ( .D(n2244), .CK(clk), .Q(n1727), .QN(n1290) );
  DFFX1 stg_reg_reg_1__30_ ( .D(n2213), .CK(clk), .Q(n1676), .QN(n1433) );
  DFFX1 stg_reg_reg_1__31_ ( .D(n2212), .CK(clk), .Q(n1679), .QN(n1426) );
  DFFX1 stg_reg_reg_12__13_ ( .D(n2134), .CK(clk), .Q(n1451), .QN(n10730) );
  DFFX1 stg_reg_reg_8__13_ ( .D(n2166), .CK(clk), .Q(n1450), .QN(n10720) );
  DFFX1 stg_reg_reg_12__14_ ( .D(n2133), .CK(clk), .Q(n1454), .QN(n10680) );
  DFFX1 stg_reg_reg_8__14_ ( .D(n2165), .CK(clk), .Q(n1453), .QN(n10670) );
  DFFX1 stg_reg_reg_12__15_ ( .D(n2132), .CK(clk), .Q(n1457), .QN(n10630) );
  DFFX1 stg_reg_reg_8__15_ ( .D(n2164), .CK(clk), .Q(n1456), .QN(n10620) );
  DFFQX1 stg_reg_reg_4__13_ ( .D(n2102), .CK(clk), .Q(stg_reg[141]) );
  DFFQX1 stg_reg_reg_4__14_ ( .D(n2101), .CK(clk), .Q(stg_reg[142]) );
  DFFQX1 stg_reg_reg_4__15_ ( .D(n2100), .CK(clk), .Q(stg_reg[143]) );
  DFFX1 stg_reg_reg_1__14_ ( .D(n2229), .CK(clk), .Q(n1500), .QN(n160) );
  DFFX1 stg_reg_reg_1__15_ ( .D(n2228), .CK(clk), .Q(n1503), .QN(n171) );
  DFFX1 stg_reg_reg_2__14_ ( .D(n2261), .CK(clk), .Q(n1548), .QN(n156) );
  DFFX1 stg_reg_reg_2__15_ ( .D(n2260), .CK(clk), .Q(n1551), .QN(n168) );
  DFFX1 stg_reg_reg_0__13_ ( .D(n2198), .CK(clk), .Q(n1449), .QN(n159) );
  DFFX1 stg_reg_reg_0__14_ ( .D(n2197), .CK(clk), .Q(n1452), .QN(n161) );
  DFFX1 stg_reg_reg_0__15_ ( .D(n2196), .CK(clk), .Q(n1455), .QN(n170) );
  DFFX1 stg_reg_reg_3__14_ ( .D(n2293), .CK(clk), .Q(n1591), .QN(n157) );
  DFFX1 stg_reg_reg_3__15_ ( .D(n2292), .CK(clk), .Q(n1593), .QN(n169) );
  DFFQX1 data_reg_0__14_ ( .D(data_1__14_), .CK(clk), .Q(data_0__14_) );
  DFFQX1 data_reg_0__13_ ( .D(data_1__13_), .CK(clk), .Q(data_0__13_) );
  DFFQX1 data_reg_0__12_ ( .D(data_1__12_), .CK(clk), .Q(data_0__12_) );
  DFFQX1 data_reg_0__11_ ( .D(data_1__11_), .CK(clk), .Q(data_0__11_) );
  DFFQX1 data_reg_0__10_ ( .D(data_1__10_), .CK(clk), .Q(data_0__10_) );
  DFFQX1 data_reg_0__9_ ( .D(data_1__9_), .CK(clk), .Q(data_0__9_) );
  DFFQX1 data_reg_0__8_ ( .D(data_1__8_), .CK(clk), .Q(data_0__8_) );
  DFFQX1 data_reg_7__15_ ( .D(data_8__15_), .CK(clk), .Q(data_7__15_) );
  DFFQX1 data_reg_6__15_ ( .D(data_7__15_), .CK(clk), .Q(data_6__15_) );
  DFFQX1 data_reg_5__15_ ( .D(data_6__15_), .CK(clk), .Q(data_5__15_) );
  DFFQX1 data_reg_4__15_ ( .D(data_5__15_), .CK(clk), .Q(data_4__15_) );
  DFFQX1 data_reg_7__14_ ( .D(data_8__14_), .CK(clk), .Q(data_7__14_) );
  DFFQX1 data_reg_6__14_ ( .D(data_7__14_), .CK(clk), .Q(data_6__14_) );
  DFFQX1 data_reg_5__14_ ( .D(data_6__14_), .CK(clk), .Q(data_5__14_) );
  DFFQX1 data_reg_4__14_ ( .D(data_5__14_), .CK(clk), .Q(data_4__14_) );
  DFFQX1 data_reg_7__13_ ( .D(data_8__13_), .CK(clk), .Q(data_7__13_) );
  DFFQX1 data_reg_6__13_ ( .D(data_7__13_), .CK(clk), .Q(data_6__13_) );
  DFFQX1 data_reg_5__13_ ( .D(data_6__13_), .CK(clk), .Q(data_5__13_) );
  DFFQX1 data_reg_4__13_ ( .D(data_5__13_), .CK(clk), .Q(data_4__13_) );
  DFFQX1 data_reg_7__12_ ( .D(data_8__12_), .CK(clk), .Q(data_7__12_) );
  DFFQX1 data_reg_6__12_ ( .D(data_7__12_), .CK(clk), .Q(data_6__12_) );
  DFFQX1 data_reg_5__12_ ( .D(data_6__12_), .CK(clk), .Q(data_5__12_) );
  DFFQX1 data_reg_4__12_ ( .D(data_5__12_), .CK(clk), .Q(data_4__12_) );
  DFFQX1 data_reg_7__11_ ( .D(data_8__11_), .CK(clk), .Q(data_7__11_) );
  DFFQX1 data_reg_6__11_ ( .D(data_7__11_), .CK(clk), .Q(data_6__11_) );
  DFFQX1 data_reg_5__11_ ( .D(data_6__11_), .CK(clk), .Q(data_5__11_) );
  DFFQX1 data_reg_4__11_ ( .D(data_5__11_), .CK(clk), .Q(data_4__11_) );
  DFFQX1 data_reg_7__10_ ( .D(data_8__10_), .CK(clk), .Q(data_7__10_) );
  DFFQX1 data_reg_6__10_ ( .D(data_7__10_), .CK(clk), .Q(data_6__10_) );
  DFFQX1 data_reg_5__10_ ( .D(data_6__10_), .CK(clk), .Q(data_5__10_) );
  DFFQX1 data_reg_4__10_ ( .D(data_5__10_), .CK(clk), .Q(data_4__10_) );
  DFFQX1 data_reg_7__9_ ( .D(data_8__9_), .CK(clk), .Q(data_7__9_) );
  DFFQX1 data_reg_6__9_ ( .D(data_7__9_), .CK(clk), .Q(data_6__9_) );
  DFFQX1 data_reg_5__9_ ( .D(data_6__9_), .CK(clk), .Q(data_5__9_) );
  DFFQX1 data_reg_4__9_ ( .D(data_5__9_), .CK(clk), .Q(data_4__9_) );
  DFFQX1 data_reg_4__8_ ( .D(data_5__8_), .CK(clk), .Q(data_4__8_) );
  DFFQX1 data_reg_3__15_ ( .D(data_4__15_), .CK(clk), .Q(data_3__15_) );
  DFFQX1 data_reg_2__15_ ( .D(data_3__15_), .CK(clk), .Q(data_2__15_) );
  DFFQX1 data_reg_1__15_ ( .D(data_2__15_), .CK(clk), .Q(data_1__15_) );
  DFFQX1 data_reg_3__14_ ( .D(data_4__14_), .CK(clk), .Q(data_3__14_) );
  DFFQX1 data_reg_2__14_ ( .D(data_3__14_), .CK(clk), .Q(data_2__14_) );
  DFFQX1 data_reg_1__14_ ( .D(data_2__14_), .CK(clk), .Q(data_1__14_) );
  DFFQX1 data_reg_3__13_ ( .D(data_4__13_), .CK(clk), .Q(data_3__13_) );
  DFFQX1 data_reg_2__13_ ( .D(data_3__13_), .CK(clk), .Q(data_2__13_) );
  DFFQX1 data_reg_1__13_ ( .D(data_2__13_), .CK(clk), .Q(data_1__13_) );
  DFFQX1 data_reg_3__12_ ( .D(data_4__12_), .CK(clk), .Q(data_3__12_) );
  DFFQX1 data_reg_2__12_ ( .D(data_3__12_), .CK(clk), .Q(data_2__12_) );
  DFFQX1 data_reg_1__12_ ( .D(data_2__12_), .CK(clk), .Q(data_1__12_) );
  DFFQX1 data_reg_3__11_ ( .D(data_4__11_), .CK(clk), .Q(data_3__11_) );
  DFFQX1 data_reg_2__11_ ( .D(data_3__11_), .CK(clk), .Q(data_2__11_) );
  DFFQX1 data_reg_1__11_ ( .D(data_2__11_), .CK(clk), .Q(data_1__11_) );
  DFFQX1 data_reg_3__10_ ( .D(data_4__10_), .CK(clk), .Q(data_3__10_) );
  DFFQX1 data_reg_2__10_ ( .D(data_3__10_), .CK(clk), .Q(data_2__10_) );
  DFFQX1 data_reg_1__10_ ( .D(data_2__10_), .CK(clk), .Q(data_1__10_) );
  DFFQX1 data_reg_3__9_ ( .D(data_4__9_), .CK(clk), .Q(data_3__9_) );
  DFFQX1 data_reg_2__9_ ( .D(data_3__9_), .CK(clk), .Q(data_2__9_) );
  DFFQX1 data_reg_1__9_ ( .D(data_2__9_), .CK(clk), .Q(data_1__9_) );
  DFFQX1 data_reg_3__8_ ( .D(data_4__8_), .CK(clk), .Q(data_3__8_) );
  DFFQX1 data_reg_2__8_ ( .D(data_3__8_), .CK(clk), .Q(data_2__8_) );
  DFFQX1 data_reg_1__8_ ( .D(data_2__8_), .CK(clk), .Q(data_1__8_) );
  DFFQX1 data_reg_11__15_ ( .D(data_12__15_), .CK(clk), .Q(data_11__15_) );
  DFFQX1 data_reg_10__15_ ( .D(data_11__15_), .CK(clk), .Q(data_10__15_) );
  DFFQX1 data_reg_9__15_ ( .D(data_10__15_), .CK(clk), .Q(data_9__15_) );
  DFFQX1 data_reg_11__14_ ( .D(data_12__14_), .CK(clk), .Q(data_11__14_) );
  DFFQX1 data_reg_10__14_ ( .D(data_11__14_), .CK(clk), .Q(data_10__14_) );
  DFFQX1 data_reg_9__14_ ( .D(data_10__14_), .CK(clk), .Q(data_9__14_) );
  DFFQX1 data_reg_8__14_ ( .D(data_9__14_), .CK(clk), .Q(data_8__14_) );
  DFFQX1 data_reg_11__13_ ( .D(data_12__13_), .CK(clk), .Q(data_11__13_) );
  DFFQX1 data_reg_10__13_ ( .D(data_11__13_), .CK(clk), .Q(data_10__13_) );
  DFFQX1 data_reg_9__13_ ( .D(data_10__13_), .CK(clk), .Q(data_9__13_) );
  DFFQX1 data_reg_8__13_ ( .D(data_9__13_), .CK(clk), .Q(data_8__13_) );
  DFFQX1 data_reg_11__12_ ( .D(data_12__12_), .CK(clk), .Q(data_11__12_) );
  DFFQX1 data_reg_10__12_ ( .D(data_11__12_), .CK(clk), .Q(data_10__12_) );
  DFFQX1 data_reg_9__12_ ( .D(data_10__12_), .CK(clk), .Q(data_9__12_) );
  DFFQX1 data_reg_8__12_ ( .D(data_9__12_), .CK(clk), .Q(data_8__12_) );
  DFFQX1 data_reg_11__11_ ( .D(data_12__11_), .CK(clk), .Q(data_11__11_) );
  DFFQX1 data_reg_10__11_ ( .D(data_11__11_), .CK(clk), .Q(data_10__11_) );
  DFFQX1 data_reg_9__11_ ( .D(data_10__11_), .CK(clk), .Q(data_9__11_) );
  DFFQX1 data_reg_8__11_ ( .D(data_9__11_), .CK(clk), .Q(data_8__11_) );
  DFFQX1 data_reg_11__10_ ( .D(data_12__10_), .CK(clk), .Q(data_11__10_) );
  DFFQX1 data_reg_10__10_ ( .D(data_11__10_), .CK(clk), .Q(data_10__10_) );
  DFFQX1 data_reg_9__10_ ( .D(data_10__10_), .CK(clk), .Q(data_9__10_) );
  DFFQX1 data_reg_8__10_ ( .D(data_9__10_), .CK(clk), .Q(data_8__10_) );
  DFFQX1 data_reg_11__9_ ( .D(data_12__9_), .CK(clk), .Q(data_11__9_) );
  DFFQX1 data_reg_10__9_ ( .D(data_11__9_), .CK(clk), .Q(data_10__9_) );
  DFFQX1 data_reg_9__9_ ( .D(data_10__9_), .CK(clk), .Q(data_9__9_) );
  DFFQX1 data_reg_8__9_ ( .D(data_9__9_), .CK(clk), .Q(data_8__9_) );
  DFFQX1 data_reg_11__8_ ( .D(data_12__8_), .CK(clk), .Q(data_11__8_) );
  DFFQX1 data_reg_10__8_ ( .D(data_11__8_), .CK(clk), .Q(data_10__8_) );
  DFFQX1 data_reg_9__8_ ( .D(data_10__8_), .CK(clk), .Q(data_9__8_) );
  DFFQX1 data_reg_8__8_ ( .D(data_9__8_), .CK(clk), .Q(data_8__8_) );
  DFFQX1 data_reg_14__15_ ( .D(fir_d[15]), .CK(clk), .Q(data_14__15_) );
  DFFQX1 data_reg_13__15_ ( .D(data_14__15_), .CK(clk), .Q(data_13__15_) );
  DFFQX1 data_reg_12__15_ ( .D(data_13__15_), .CK(clk), .Q(data_12__15_) );
  DFFQX1 data_reg_14__14_ ( .D(fir_d[14]), .CK(clk), .Q(data_14__14_) );
  DFFQX1 data_reg_13__14_ ( .D(data_14__14_), .CK(clk), .Q(data_13__14_) );
  DFFQX1 data_reg_12__14_ ( .D(data_13__14_), .CK(clk), .Q(data_12__14_) );
  DFFQX1 data_reg_14__13_ ( .D(fir_d[13]), .CK(clk), .Q(data_14__13_) );
  DFFQX1 data_reg_13__13_ ( .D(data_14__13_), .CK(clk), .Q(data_13__13_) );
  DFFQX1 data_reg_12__13_ ( .D(data_13__13_), .CK(clk), .Q(data_12__13_) );
  DFFQX1 data_reg_14__12_ ( .D(fir_d[12]), .CK(clk), .Q(data_14__12_) );
  DFFQX1 data_reg_13__12_ ( .D(data_14__12_), .CK(clk), .Q(data_13__12_) );
  DFFQX1 data_reg_12__12_ ( .D(data_13__12_), .CK(clk), .Q(data_12__12_) );
  DFFQX1 data_reg_14__11_ ( .D(fir_d[11]), .CK(clk), .Q(data_14__11_) );
  DFFQX1 data_reg_13__11_ ( .D(data_14__11_), .CK(clk), .Q(data_13__11_) );
  DFFQX1 data_reg_12__11_ ( .D(data_13__11_), .CK(clk), .Q(data_12__11_) );
  DFFQX1 data_reg_14__10_ ( .D(fir_d[10]), .CK(clk), .Q(data_14__10_) );
  DFFQX1 data_reg_13__10_ ( .D(data_14__10_), .CK(clk), .Q(data_13__10_) );
  DFFQX1 data_reg_12__10_ ( .D(data_13__10_), .CK(clk), .Q(data_12__10_) );
  DFFQX1 data_reg_14__9_ ( .D(fir_d[9]), .CK(clk), .Q(data_14__9_) );
  DFFQX1 data_reg_13__9_ ( .D(data_14__9_), .CK(clk), .Q(data_13__9_) );
  DFFQX1 data_reg_12__9_ ( .D(data_13__9_), .CK(clk), .Q(data_12__9_) );
  DFFQX1 data_reg_12__8_ ( .D(data_13__8_), .CK(clk), .Q(data_12__8_) );
  DFFQX1 stg_reg_reg_4__21_ ( .D(n3219), .CK(clk), .Q(stg_reg[149]) );
  DFFQX1 stg_reg_reg_4__22_ ( .D(n3218), .CK(clk), .Q(stg_reg[150]) );
  DFFQX1 stg_reg_reg_4__23_ ( .D(n3217), .CK(clk), .Q(stg_reg[151]) );
  DFFQX1 stg_reg_reg_4__24_ ( .D(n3216), .CK(clk), .Q(stg_reg[152]) );
  DFFQX1 stg_reg_reg_4__25_ ( .D(n3215), .CK(clk), .Q(stg_reg[153]) );
  DFFQX1 stg_reg_reg_4__26_ ( .D(n3214), .CK(clk), .Q(stg_reg[154]) );
  DFFQX1 stg_reg_reg_4__27_ ( .D(n3213), .CK(clk), .Q(stg_reg[155]) );
  DFFX1 stg_reg_reg_3__22_ ( .D(n2285), .CK(clk), .Q(n1781), .QN(n2639) );
  DFFX1 stg_reg_reg_3__23_ ( .D(n2284), .CK(clk), .Q(n1783), .QN(n2630) );
  DFFX1 stg_reg_reg_3__24_ ( .D(n2283), .CK(clk), .Q(n1785), .QN(n2621) );
  DFFX1 stg_reg_reg_3__25_ ( .D(n2282), .CK(clk), .Q(n1787), .QN(n2612) );
  DFFX1 stg_reg_reg_3__26_ ( .D(n2281), .CK(clk), .Q(n1759), .QN(n2603) );
  DFFX1 stg_reg_reg_3__27_ ( .D(n2280), .CK(clk), .Q(n1761), .QN(n2594) );
  DFFX1 stg_reg_reg_3__28_ ( .D(n2279), .CK(clk), .Q(n1763), .QN(n2585) );
  DFFX1 stg_reg_reg_3__29_ ( .D(n2278), .CK(clk), .Q(n1765), .QN(n2576) );
  DFFX1 stg_reg_reg_12__21_ ( .D(n2126), .CK(clk), .Q(n1648), .QN(n1238) );
  DFFX1 stg_reg_reg_8__21_ ( .D(n2158), .CK(clk), .Q(n1647), .QN(n1237) );
  DFFX1 stg_reg_reg_0__21_ ( .D(n2190), .CK(clk), .Q(n1646), .QN(n1234) );
  DFFX1 stg_reg_reg_12__22_ ( .D(n2125), .CK(clk), .Q(n1651), .QN(n1229) );
  DFFX1 stg_reg_reg_8__22_ ( .D(n2157), .CK(clk), .Q(n1650), .QN(n1228) );
  DFFX1 stg_reg_reg_0__22_ ( .D(n2189), .CK(clk), .Q(n1649), .QN(n1225) );
  DFFX1 stg_reg_reg_12__23_ ( .D(n2124), .CK(clk), .Q(n1654), .QN(n1220) );
  DFFX1 stg_reg_reg_8__23_ ( .D(n2156), .CK(clk), .Q(n1653), .QN(n1219) );
  DFFX1 stg_reg_reg_0__23_ ( .D(n2188), .CK(clk), .Q(n1652), .QN(n1216) );
  DFFX1 stg_reg_reg_12__24_ ( .D(n2123), .CK(clk), .Q(n1657), .QN(n1211) );
  DFFX1 stg_reg_reg_8__24_ ( .D(n2155), .CK(clk), .Q(n1656), .QN(n1210) );
  DFFX1 stg_reg_reg_0__24_ ( .D(n2187), .CK(clk), .Q(n1655), .QN(n1207) );
  DFFX1 stg_reg_reg_12__25_ ( .D(n2122), .CK(clk), .Q(n1660), .QN(n1202) );
  DFFX1 stg_reg_reg_8__25_ ( .D(n2154), .CK(clk), .Q(n1659), .QN(n1201) );
  DFFX1 stg_reg_reg_0__25_ ( .D(n2186), .CK(clk), .Q(n1658), .QN(n1198) );
  DFFX1 stg_reg_reg_12__26_ ( .D(n2121), .CK(clk), .Q(n1618), .QN(n1193) );
  DFFX1 stg_reg_reg_8__26_ ( .D(n2153), .CK(clk), .Q(n1617), .QN(n1192) );
  DFFX1 stg_reg_reg_0__26_ ( .D(n2185), .CK(clk), .Q(n1616), .QN(n1189) );
  DFFX1 stg_reg_reg_12__27_ ( .D(n2120), .CK(clk), .Q(n1621), .QN(n1184) );
  DFFX1 stg_reg_reg_8__27_ ( .D(n2152), .CK(clk), .Q(n1620), .QN(n1183) );
  DFFX1 stg_reg_reg_0__27_ ( .D(n2184), .CK(clk), .Q(n1619), .QN(n1180) );
  DFFX1 stg_reg_reg_8__28_ ( .D(n2151), .CK(clk), .Q(n1623), .QN(n1174) );
  DFFX1 stg_reg_reg_0__28_ ( .D(n2183), .CK(clk), .Q(n1622), .QN(n1171) );
  DFFX1 stg_reg_reg_2__22_ ( .D(n2253), .CK(clk), .Q(n1745), .QN(n1366) );
  DFFX1 stg_reg_reg_2__23_ ( .D(n2252), .CK(clk), .Q(n1748), .QN(n1358) );
  DFFX1 stg_reg_reg_2__24_ ( .D(n2251), .CK(clk), .Q(n1751), .QN(n1350) );
  DFFX1 stg_reg_reg_2__25_ ( .D(n2250), .CK(clk), .Q(n1754), .QN(n1341) );
  DFFX1 stg_reg_reg_2__26_ ( .D(n2249), .CK(clk), .Q(n1712), .QN(n1332) );
  DFFX1 stg_reg_reg_2__27_ ( .D(n2248), .CK(clk), .Q(n1715), .QN(n1323) );
  DFFX1 stg_reg_reg_2__28_ ( .D(n2247), .CK(clk), .Q(n1718), .QN(n1314) );
  DFFX1 stg_reg_reg_2__29_ ( .D(n2246), .CK(clk), .Q(n1721), .QN(n1305) );
  DFFX1 stg_reg_reg_1__22_ ( .D(n2221), .CK(clk), .Q(n1697), .QN(n2343) );
  DFFX1 stg_reg_reg_1__23_ ( .D(n2220), .CK(clk), .Q(n1700), .QN(n2336) );
  DFFX1 stg_reg_reg_1__24_ ( .D(n2219), .CK(clk), .Q(n1703), .QN(n2329) );
  DFFX1 stg_reg_reg_1__25_ ( .D(n2218), .CK(clk), .Q(n1706), .QN(n2322) );
  DFFX1 stg_reg_reg_1__26_ ( .D(n2217), .CK(clk), .Q(n1664), .QN(n2315) );
  DFFX1 stg_reg_reg_1__27_ ( .D(n2216), .CK(clk), .Q(n1667), .QN(n1812) );
  DFFX1 stg_reg_reg_1__28_ ( .D(n2215), .CK(clk), .Q(n1670), .QN(n1803) );
  DFFX1 stg_reg_reg_1__29_ ( .D(n2214), .CK(clk), .Q(n1673), .QN(n1796) );
  DFFX1 stg_reg_reg_12__5_ ( .D(n2142), .CK(clk), .Q(n1472), .QN(n11170) );
  DFFX1 stg_reg_reg_8__5_ ( .D(n2174), .CK(clk), .Q(n1471), .QN(n11160) );
  DFFX1 stg_reg_reg_12__6_ ( .D(n2141), .CK(clk), .Q(n1475), .QN(n11110) );
  DFFX1 stg_reg_reg_8__6_ ( .D(n2173), .CK(clk), .Q(n1474), .QN(n11100) );
  DFFX1 stg_reg_reg_12__7_ ( .D(n2140), .CK(clk), .Q(n1478), .QN(n11050) );
  DFFX1 stg_reg_reg_8__7_ ( .D(n2172), .CK(clk), .Q(n1477), .QN(n11040) );
  DFFX1 stg_reg_reg_12__8_ ( .D(n2139), .CK(clk), .Q(n1481), .QN(n10990) );
  DFFX1 stg_reg_reg_8__8_ ( .D(n2171), .CK(clk), .Q(n1480), .QN(n10980) );
  DFFX1 stg_reg_reg_12__9_ ( .D(n2138), .CK(clk), .Q(n1484), .QN(n10930) );
  DFFX1 stg_reg_reg_8__9_ ( .D(n2170), .CK(clk), .Q(n1483), .QN(n10920) );
  DFFX1 stg_reg_reg_12__10_ ( .D(n2137), .CK(clk), .Q(n1442), .QN(n10880) );
  DFFX1 stg_reg_reg_8__10_ ( .D(n2169), .CK(clk), .Q(n1441), .QN(n10870) );
  DFFX1 stg_reg_reg_12__11_ ( .D(n2136), .CK(clk), .Q(n1445), .QN(n10830) );
  DFFX1 stg_reg_reg_8__11_ ( .D(n2168), .CK(clk), .Q(n1444), .QN(n10820) );
  DFFX1 stg_reg_reg_12__12_ ( .D(n2135), .CK(clk), .Q(n1448), .QN(n10780) );
  DFFX1 stg_reg_reg_8__12_ ( .D(n2167), .CK(clk), .Q(n1447), .QN(n10770) );
  DFFQX1 stg_reg_reg_4__5_ ( .D(n2110), .CK(clk), .Q(stg_reg[133]) );
  DFFQX1 stg_reg_reg_4__6_ ( .D(n2109), .CK(clk), .Q(stg_reg[134]) );
  DFFQX1 stg_reg_reg_4__7_ ( .D(n2108), .CK(clk), .Q(stg_reg[135]) );
  DFFQX1 stg_reg_reg_4__8_ ( .D(n2107), .CK(clk), .Q(stg_reg[136]) );
  DFFQX1 stg_reg_reg_4__9_ ( .D(n2106), .CK(clk), .Q(stg_reg[137]) );
  DFFQX1 stg_reg_reg_4__10_ ( .D(n2105), .CK(clk), .Q(stg_reg[138]) );
  DFFQX1 stg_reg_reg_4__11_ ( .D(n2104), .CK(clk), .Q(stg_reg[139]) );
  DFFQX1 stg_reg_reg_4__12_ ( .D(n2103), .CK(clk), .Q(stg_reg[140]) );
  DFFX1 stg_reg_reg_1__6_ ( .D(n2237), .CK(clk), .Q(n1521), .QN(n2429) );
  DFFX1 stg_reg_reg_1__7_ ( .D(n2236), .CK(clk), .Q(n1524), .QN(n2424) );
  DFFX1 stg_reg_reg_1__8_ ( .D(n2235), .CK(clk), .Q(n1527), .QN(n2419) );
  DFFX1 stg_reg_reg_1__9_ ( .D(n2234), .CK(clk), .Q(n1530), .QN(n141) );
  DFFX1 stg_reg_reg_1__10_ ( .D(n2233), .CK(clk), .Q(n1488), .QN(n142) );
  DFFX1 stg_reg_reg_1__11_ ( .D(n2232), .CK(clk), .Q(n1491), .QN(n143) );
  DFFX1 stg_reg_reg_1__12_ ( .D(n2231), .CK(clk), .Q(n1494), .QN(n144) );
  DFFX1 stg_reg_reg_1__13_ ( .D(n2230), .CK(clk), .Q(n1497), .QN(n158) );
  DFFX1 stg_reg_reg_2__6_ ( .D(n2269), .CK(clk), .Q(n1569), .QN(n3116) );
  DFFX1 stg_reg_reg_2__7_ ( .D(n2268), .CK(clk), .Q(n1572), .QN(n3112) );
  DFFX1 stg_reg_reg_2__8_ ( .D(n2267), .CK(clk), .Q(n1575), .QN(n3107) );
  DFFX1 stg_reg_reg_2__9_ ( .D(n2266), .CK(clk), .Q(n1578), .QN(n127) );
  DFFX1 stg_reg_reg_2__10_ ( .D(n2265), .CK(clk), .Q(n1536), .QN(n133) );
  DFFX1 stg_reg_reg_2__11_ ( .D(n2264), .CK(clk), .Q(n1539), .QN(n135) );
  DFFX1 stg_reg_reg_2__12_ ( .D(n2263), .CK(clk), .Q(n1542), .QN(n137) );
  DFFX1 stg_reg_reg_2__13_ ( .D(n2262), .CK(clk), .Q(n1545), .QN(n154) );
  DFFX1 stg_reg_reg_0__5_ ( .D(n2206), .CK(clk), .Q(n1470), .QN(n11130) );
  DFFX1 stg_reg_reg_0__6_ ( .D(n2205), .CK(clk), .Q(n1473), .QN(n11070) );
  DFFX1 stg_reg_reg_0__7_ ( .D(n2204), .CK(clk), .Q(n1476), .QN(n11010) );
  DFFX1 stg_reg_reg_0__8_ ( .D(n2203), .CK(clk), .Q(n1479), .QN(n10950) );
  DFFX1 stg_reg_reg_0__9_ ( .D(n2202), .CK(clk), .Q(n1482), .QN(n139) );
  DFFX1 stg_reg_reg_0__10_ ( .D(n2201), .CK(clk), .Q(n1440), .QN(n140) );
  DFFX1 stg_reg_reg_0__11_ ( .D(n2200), .CK(clk), .Q(n1443), .QN(n145) );
  DFFX1 stg_reg_reg_0__12_ ( .D(n2199), .CK(clk), .Q(n1446), .QN(n146) );
  DFFX1 stg_reg_reg_3__6_ ( .D(n2301), .CK(clk), .Q(n1605), .QN(n2515) );
  DFFX1 stg_reg_reg_3__7_ ( .D(n2300), .CK(clk), .Q(n1607), .QN(n2509) );
  DFFX1 stg_reg_reg_3__8_ ( .D(n2299), .CK(clk), .Q(n1609), .QN(n2503) );
  DFFX1 stg_reg_reg_3__9_ ( .D(n2298), .CK(clk), .Q(n1611), .QN(n128) );
  DFFX1 stg_reg_reg_3__10_ ( .D(n2297), .CK(clk), .Q(n1583), .QN(n134) );
  DFFX1 stg_reg_reg_3__11_ ( .D(n2296), .CK(clk), .Q(n1585), .QN(n136) );
  DFFX1 stg_reg_reg_3__12_ ( .D(n2295), .CK(clk), .Q(n1587), .QN(n138) );
  DFFX1 stg_reg_reg_3__13_ ( .D(n2294), .CK(clk), .Q(n1589), .QN(n155) );
  DFFQX1 data_reg_0__7_ ( .D(data_1__7_), .CK(clk), .Q(data_0__7_) );
  DFFQX1 data_reg_0__6_ ( .D(data_1__6_), .CK(clk), .Q(data_0__6_) );
  DFFQX1 data_reg_0__5_ ( .D(data_1__5_), .CK(clk), .Q(data_0__5_) );
  DFFQX1 data_reg_0__4_ ( .D(data_1__4_), .CK(clk), .Q(data_0__4_) );
  DFFQX1 data_reg_0__3_ ( .D(data_1__3_), .CK(clk), .Q(data_0__3_) );
  DFFQX1 data_reg_0__2_ ( .D(data_1__2_), .CK(clk), .Q(data_0__2_) );
  DFFQX1 data_reg_0__1_ ( .D(data_1__1_), .CK(clk), .Q(data_0__1_) );
  DFFQX1 data_reg_7__8_ ( .D(data_8__8_), .CK(clk), .Q(data_7__8_) );
  DFFQX1 data_reg_6__8_ ( .D(data_7__8_), .CK(clk), .Q(data_6__8_) );
  DFFQX1 data_reg_5__8_ ( .D(data_6__8_), .CK(clk), .Q(data_5__8_) );
  DFFQX1 data_reg_7__7_ ( .D(data_8__7_), .CK(clk), .Q(data_7__7_) );
  DFFQX1 data_reg_6__7_ ( .D(data_7__7_), .CK(clk), .Q(data_6__7_) );
  DFFQX1 data_reg_5__7_ ( .D(data_6__7_), .CK(clk), .Q(data_5__7_) );
  DFFQX1 data_reg_4__7_ ( .D(data_5__7_), .CK(clk), .Q(data_4__7_) );
  DFFQX1 data_reg_7__6_ ( .D(data_8__6_), .CK(clk), .Q(data_7__6_) );
  DFFQX1 data_reg_6__6_ ( .D(data_7__6_), .CK(clk), .Q(data_6__6_) );
  DFFQX1 data_reg_5__6_ ( .D(data_6__6_), .CK(clk), .Q(data_5__6_) );
  DFFQX1 data_reg_4__6_ ( .D(data_5__6_), .CK(clk), .Q(data_4__6_) );
  DFFQX1 data_reg_7__5_ ( .D(data_8__5_), .CK(clk), .Q(data_7__5_) );
  DFFQX1 data_reg_6__5_ ( .D(data_7__5_), .CK(clk), .Q(data_6__5_) );
  DFFQX1 data_reg_5__5_ ( .D(data_6__5_), .CK(clk), .Q(data_5__5_) );
  DFFQX1 data_reg_4__5_ ( .D(data_5__5_), .CK(clk), .Q(data_4__5_) );
  DFFQX1 data_reg_7__4_ ( .D(data_8__4_), .CK(clk), .Q(data_7__4_) );
  DFFQX1 data_reg_6__4_ ( .D(data_7__4_), .CK(clk), .Q(data_6__4_) );
  DFFQX1 data_reg_5__4_ ( .D(data_6__4_), .CK(clk), .Q(data_5__4_) );
  DFFQX1 data_reg_4__4_ ( .D(data_5__4_), .CK(clk), .Q(data_4__4_) );
  DFFQX1 data_reg_7__3_ ( .D(data_8__3_), .CK(clk), .Q(data_7__3_) );
  DFFQX1 data_reg_6__3_ ( .D(data_7__3_), .CK(clk), .Q(data_6__3_) );
  DFFQX1 data_reg_5__3_ ( .D(data_6__3_), .CK(clk), .Q(data_5__3_) );
  DFFQX1 data_reg_4__3_ ( .D(data_5__3_), .CK(clk), .Q(data_4__3_) );
  DFFQX1 data_reg_7__2_ ( .D(data_8__2_), .CK(clk), .Q(data_7__2_) );
  DFFQX1 data_reg_6__2_ ( .D(data_7__2_), .CK(clk), .Q(data_6__2_) );
  DFFQX1 data_reg_5__2_ ( .D(data_6__2_), .CK(clk), .Q(data_5__2_) );
  DFFQX1 data_reg_4__2_ ( .D(data_5__2_), .CK(clk), .Q(data_4__2_) );
  DFFQX1 data_reg_7__1_ ( .D(data_8__1_), .CK(clk), .Q(data_7__1_) );
  DFFQX1 data_reg_6__1_ ( .D(data_7__1_), .CK(clk), .Q(data_6__1_) );
  DFFQX1 data_reg_5__1_ ( .D(data_6__1_), .CK(clk), .Q(data_5__1_) );
  DFFQX1 data_reg_4__1_ ( .D(data_5__1_), .CK(clk), .Q(data_4__1_) );
  DFFQX1 data_reg_3__7_ ( .D(data_4__7_), .CK(clk), .Q(data_3__7_) );
  DFFQX1 data_reg_2__7_ ( .D(data_3__7_), .CK(clk), .Q(data_2__7_) );
  DFFQX1 data_reg_1__7_ ( .D(data_2__7_), .CK(clk), .Q(data_1__7_) );
  DFFQX1 data_reg_3__6_ ( .D(data_4__6_), .CK(clk), .Q(data_3__6_) );
  DFFQX1 data_reg_2__6_ ( .D(data_3__6_), .CK(clk), .Q(data_2__6_) );
  DFFQX1 data_reg_1__6_ ( .D(data_2__6_), .CK(clk), .Q(data_1__6_) );
  DFFQX1 data_reg_3__5_ ( .D(data_4__5_), .CK(clk), .Q(data_3__5_) );
  DFFQX1 data_reg_2__5_ ( .D(data_3__5_), .CK(clk), .Q(data_2__5_) );
  DFFQX1 data_reg_1__5_ ( .D(data_2__5_), .CK(clk), .Q(data_1__5_) );
  DFFQX1 data_reg_3__4_ ( .D(data_4__4_), .CK(clk), .Q(data_3__4_) );
  DFFQX1 data_reg_2__4_ ( .D(data_3__4_), .CK(clk), .Q(data_2__4_) );
  DFFQX1 data_reg_1__4_ ( .D(data_2__4_), .CK(clk), .Q(data_1__4_) );
  DFFQX1 data_reg_3__3_ ( .D(data_4__3_), .CK(clk), .Q(data_3__3_) );
  DFFQX1 data_reg_2__3_ ( .D(data_3__3_), .CK(clk), .Q(data_2__3_) );
  DFFQX1 data_reg_1__3_ ( .D(data_2__3_), .CK(clk), .Q(data_1__3_) );
  DFFQX1 data_reg_3__2_ ( .D(data_4__2_), .CK(clk), .Q(data_3__2_) );
  DFFQX1 data_reg_2__2_ ( .D(data_3__2_), .CK(clk), .Q(data_2__2_) );
  DFFQX1 data_reg_1__2_ ( .D(data_2__2_), .CK(clk), .Q(data_1__2_) );
  DFFQX1 data_reg_3__1_ ( .D(data_4__1_), .CK(clk), .Q(data_3__1_) );
  DFFQX1 data_reg_2__1_ ( .D(data_3__1_), .CK(clk), .Q(data_2__1_) );
  DFFQX1 data_reg_1__1_ ( .D(data_2__1_), .CK(clk), .Q(data_1__1_) );
  DFFQX1 data_reg_11__0_ ( .D(data_12__0_), .CK(clk), .Q(data_11__0_) );
  DFFQX1 data_reg_10__0_ ( .D(data_11__0_), .CK(clk), .Q(data_10__0_) );
  DFFQX1 data_reg_9__0_ ( .D(data_10__0_), .CK(clk), .Q(data_9__0_) );
  DFFQX1 data_reg_8__0_ ( .D(data_9__0_), .CK(clk), .Q(data_8__0_) );
  DFFQX1 data_reg_11__7_ ( .D(data_12__7_), .CK(clk), .Q(data_11__7_) );
  DFFQX1 data_reg_10__7_ ( .D(data_11__7_), .CK(clk), .Q(data_10__7_) );
  DFFQX1 data_reg_9__7_ ( .D(data_10__7_), .CK(clk), .Q(data_9__7_) );
  DFFQX1 data_reg_8__7_ ( .D(data_9__7_), .CK(clk), .Q(data_8__7_) );
  DFFQX1 data_reg_11__6_ ( .D(data_12__6_), .CK(clk), .Q(data_11__6_) );
  DFFQX1 data_reg_10__6_ ( .D(data_11__6_), .CK(clk), .Q(data_10__6_) );
  DFFQX1 data_reg_9__6_ ( .D(data_10__6_), .CK(clk), .Q(data_9__6_) );
  DFFQX1 data_reg_8__6_ ( .D(data_9__6_), .CK(clk), .Q(data_8__6_) );
  DFFQX1 data_reg_11__5_ ( .D(data_12__5_), .CK(clk), .Q(data_11__5_) );
  DFFQX1 data_reg_10__5_ ( .D(data_11__5_), .CK(clk), .Q(data_10__5_) );
  DFFQX1 data_reg_9__5_ ( .D(data_10__5_), .CK(clk), .Q(data_9__5_) );
  DFFQX1 data_reg_8__5_ ( .D(data_9__5_), .CK(clk), .Q(data_8__5_) );
  DFFQX1 data_reg_11__4_ ( .D(data_12__4_), .CK(clk), .Q(data_11__4_) );
  DFFQX1 data_reg_10__4_ ( .D(data_11__4_), .CK(clk), .Q(data_10__4_) );
  DFFQX1 data_reg_9__4_ ( .D(data_10__4_), .CK(clk), .Q(data_9__4_) );
  DFFQX1 data_reg_8__4_ ( .D(data_9__4_), .CK(clk), .Q(data_8__4_) );
  DFFQX1 data_reg_11__3_ ( .D(data_12__3_), .CK(clk), .Q(data_11__3_) );
  DFFQX1 data_reg_10__3_ ( .D(data_11__3_), .CK(clk), .Q(data_10__3_) );
  DFFQX1 data_reg_9__3_ ( .D(data_10__3_), .CK(clk), .Q(data_9__3_) );
  DFFQX1 data_reg_8__3_ ( .D(data_9__3_), .CK(clk), .Q(data_8__3_) );
  DFFQX1 data_reg_11__2_ ( .D(data_12__2_), .CK(clk), .Q(data_11__2_) );
  DFFQX1 data_reg_10__2_ ( .D(data_11__2_), .CK(clk), .Q(data_10__2_) );
  DFFQX1 data_reg_9__2_ ( .D(data_10__2_), .CK(clk), .Q(data_9__2_) );
  DFFQX1 data_reg_8__2_ ( .D(data_9__2_), .CK(clk), .Q(data_8__2_) );
  DFFQX1 data_reg_11__1_ ( .D(data_12__1_), .CK(clk), .Q(data_11__1_) );
  DFFQX1 data_reg_10__1_ ( .D(data_11__1_), .CK(clk), .Q(data_10__1_) );
  DFFQX1 data_reg_9__1_ ( .D(data_10__1_), .CK(clk), .Q(data_9__1_) );
  DFFQX1 data_reg_8__1_ ( .D(data_9__1_), .CK(clk), .Q(data_8__1_) );
  DFFQX1 data_reg_6__0_ ( .D(data_7__0_), .CK(clk), .Q(data_6__0_) );
  DFFQX1 data_reg_5__0_ ( .D(data_6__0_), .CK(clk), .Q(data_5__0_) );
  DFFQX1 data_reg_4__0_ ( .D(data_5__0_), .CK(clk), .Q(data_4__0_) );
  DFFQX1 data_reg_14__8_ ( .D(fir_d[8]), .CK(clk), .Q(data_14__8_) );
  DFFQX1 data_reg_13__8_ ( .D(data_14__8_), .CK(clk), .Q(data_13__8_) );
  DFFQX1 data_reg_14__7_ ( .D(fir_d[7]), .CK(clk), .Q(data_14__7_) );
  DFFQX1 data_reg_13__7_ ( .D(data_14__7_), .CK(clk), .Q(data_13__7_) );
  DFFQX1 data_reg_12__7_ ( .D(data_13__7_), .CK(clk), .Q(data_12__7_) );
  DFFQX1 data_reg_14__6_ ( .D(fir_d[6]), .CK(clk), .Q(data_14__6_) );
  DFFQX1 data_reg_13__6_ ( .D(data_14__6_), .CK(clk), .Q(data_13__6_) );
  DFFQX1 data_reg_12__6_ ( .D(data_13__6_), .CK(clk), .Q(data_12__6_) );
  DFFQX1 data_reg_14__5_ ( .D(fir_d[5]), .CK(clk), .Q(data_14__5_) );
  DFFQX1 data_reg_13__5_ ( .D(data_14__5_), .CK(clk), .Q(data_13__5_) );
  DFFQX1 data_reg_12__5_ ( .D(data_13__5_), .CK(clk), .Q(data_12__5_) );
  DFFQX1 data_reg_14__4_ ( .D(fir_d[4]), .CK(clk), .Q(data_14__4_) );
  DFFQX1 data_reg_13__4_ ( .D(data_14__4_), .CK(clk), .Q(data_13__4_) );
  DFFQX1 data_reg_12__4_ ( .D(data_13__4_), .CK(clk), .Q(data_12__4_) );
  DFFQX1 data_reg_14__3_ ( .D(fir_d[3]), .CK(clk), .Q(data_14__3_) );
  DFFQX1 data_reg_13__3_ ( .D(data_14__3_), .CK(clk), .Q(data_13__3_) );
  DFFQX1 data_reg_12__3_ ( .D(data_13__3_), .CK(clk), .Q(data_12__3_) );
  DFFQX1 data_reg_14__2_ ( .D(fir_d[2]), .CK(clk), .Q(data_14__2_) );
  DFFQX1 data_reg_13__2_ ( .D(data_14__2_), .CK(clk), .Q(data_13__2_) );
  DFFQX1 data_reg_12__2_ ( .D(data_13__2_), .CK(clk), .Q(data_12__2_) );
  DFFQX1 data_reg_14__1_ ( .D(fir_d[1]), .CK(clk), .Q(data_14__1_) );
  DFFQX1 data_reg_13__1_ ( .D(data_14__1_), .CK(clk), .Q(data_13__1_) );
  DFFQX1 data_reg_12__1_ ( .D(data_13__1_), .CK(clk), .Q(data_12__1_) );
  DFFQX1 data_reg_0__0_ ( .D(data_1__0_), .CK(clk), .Q(data_0__0_) );
  DFFQX1 stg_reg_reg_4__16_ ( .D(n3224), .CK(clk), .Q(stg_reg[144]) );
  DFFQX1 stg_reg_reg_4__17_ ( .D(n3223), .CK(clk), .Q(stg_reg[145]) );
  DFFQX1 stg_reg_reg_4__18_ ( .D(n3222), .CK(clk), .Q(stg_reg[146]) );
  DFFQX1 stg_reg_reg_4__19_ ( .D(n3221), .CK(clk), .Q(stg_reg[147]) );
  DFFQX1 stg_reg_reg_4__20_ ( .D(n3220), .CK(clk), .Q(stg_reg[148]) );
  DFFX1 stg_reg_reg_3__16_ ( .D(n2291), .CK(clk), .Q(n1757), .QN(n2695) );
  DFFX1 stg_reg_reg_3__17_ ( .D(n2290), .CK(clk), .Q(n1771), .QN(n2684) );
  DFFX1 stg_reg_reg_3__18_ ( .D(n2289), .CK(clk), .Q(n1773), .QN(n2675) );
  DFFX1 stg_reg_reg_3__19_ ( .D(n2288), .CK(clk), .Q(n1775), .QN(n2666) );
  DFFX1 stg_reg_reg_3__20_ ( .D(n2287), .CK(clk), .Q(n1777), .QN(n2657) );
  DFFX1 stg_reg_reg_3__21_ ( .D(n2286), .CK(clk), .Q(n1779), .QN(n2648) );
  DFFX1 stg_reg_reg_12__16_ ( .D(n2131), .CK(clk), .Q(n1615), .QN(n1283) );
  DFFX1 stg_reg_reg_8__16_ ( .D(n2163), .CK(clk), .Q(n1614), .QN(n1282) );
  DFFX1 stg_reg_reg_0__16_ ( .D(n2195), .CK(clk), .Q(n1613), .QN(n1279) );
  DFFX1 stg_reg_reg_12__17_ ( .D(n2130), .CK(clk), .Q(n1636), .QN(n1274) );
  DFFX1 stg_reg_reg_8__17_ ( .D(n2162), .CK(clk), .Q(n1635), .QN(n1273) );
  DFFX1 stg_reg_reg_0__17_ ( .D(n2194), .CK(clk), .Q(n1634), .QN(n1270) );
  DFFX1 stg_reg_reg_12__18_ ( .D(n2129), .CK(clk), .Q(n1639), .QN(n1265) );
  DFFX1 stg_reg_reg_8__18_ ( .D(n2161), .CK(clk), .Q(n1638), .QN(n1264) );
  DFFX1 stg_reg_reg_0__18_ ( .D(n2193), .CK(clk), .Q(n1637), .QN(n1261) );
  DFFX1 stg_reg_reg_12__19_ ( .D(n2128), .CK(clk), .Q(n1642), .QN(n1256) );
  DFFX1 stg_reg_reg_8__19_ ( .D(n2160), .CK(clk), .Q(n1641), .QN(n1255) );
  DFFX1 stg_reg_reg_0__19_ ( .D(n2192), .CK(clk), .Q(n1640), .QN(n1252) );
  DFFX1 stg_reg_reg_12__20_ ( .D(n2127), .CK(clk), .Q(n1645), .QN(n1247) );
  DFFX1 stg_reg_reg_8__20_ ( .D(n2159), .CK(clk), .Q(n1644), .QN(n1246) );
  DFFX1 stg_reg_reg_0__20_ ( .D(n2191), .CK(clk), .Q(n1643), .QN(n1243) );
  DFFX1 stg_reg_reg_2__16_ ( .D(n2259), .CK(clk), .Q(n1709), .QN(n1414) );
  DFFX1 stg_reg_reg_2__17_ ( .D(n2258), .CK(clk), .Q(n1730), .QN(n1406) );
  DFFX1 stg_reg_reg_2__18_ ( .D(n2257), .CK(clk), .Q(n1733), .QN(n1398) );
  DFFX1 stg_reg_reg_2__19_ ( .D(n2256), .CK(clk), .Q(n1736), .QN(n1390) );
  DFFX1 stg_reg_reg_2__20_ ( .D(n2255), .CK(clk), .Q(n1739), .QN(n1382) );
  DFFX1 stg_reg_reg_2__21_ ( .D(n2254), .CK(clk), .Q(n1742), .QN(n1374) );
  DFFX1 stg_reg_reg_1__16_ ( .D(n2227), .CK(clk), .Q(n1661), .QN(n2385) );
  DFFX1 stg_reg_reg_1__17_ ( .D(n2226), .CK(clk), .Q(n1682), .QN(n2378) );
  DFFX1 stg_reg_reg_1__18_ ( .D(n2225), .CK(clk), .Q(n1685), .QN(n2371) );
  DFFX1 stg_reg_reg_1__19_ ( .D(n2224), .CK(clk), .Q(n1688), .QN(n2364) );
  DFFX1 stg_reg_reg_1__20_ ( .D(n2223), .CK(clk), .Q(n1691), .QN(n2357) );
  DFFX1 stg_reg_reg_1__21_ ( .D(n2222), .CK(clk), .Q(n1694), .QN(n2350) );
  DFFX1 stg_reg_reg_12__0_ ( .D(n2147), .CK(clk), .Q(n1439), .QN(n1147) );
  DFFX1 stg_reg_reg_8__0_ ( .D(n2179), .CK(clk), .Q(n1438), .QN(n1146) );
  DFFX1 stg_reg_reg_12__1_ ( .D(n2146), .CK(clk), .Q(n1460), .QN(n11410) );
  DFFX1 stg_reg_reg_8__1_ ( .D(n2178), .CK(clk), .Q(n1459), .QN(n11400) );
  DFFX1 stg_reg_reg_12__2_ ( .D(n2145), .CK(clk), .Q(n1463), .QN(n11350) );
  DFFX1 stg_reg_reg_8__2_ ( .D(n2177), .CK(clk), .Q(n1462), .QN(n11340) );
  DFFX1 stg_reg_reg_12__3_ ( .D(n2144), .CK(clk), .Q(n1466), .QN(n11290) );
  DFFX1 stg_reg_reg_8__3_ ( .D(n2176), .CK(clk), .Q(n1465), .QN(n11280) );
  DFFX1 stg_reg_reg_12__4_ ( .D(n2143), .CK(clk), .Q(n1469), .QN(n11230) );
  DFFX1 stg_reg_reg_8__4_ ( .D(n2175), .CK(clk), .Q(n1468), .QN(n11220) );
  DFFQX1 stg_reg_reg_4__0_ ( .D(n2115), .CK(clk), .Q(stg_reg[128]) );
  DFFQX1 stg_reg_reg_4__1_ ( .D(n2114), .CK(clk), .Q(stg_reg[129]) );
  DFFQX1 stg_reg_reg_4__2_ ( .D(n2113), .CK(clk), .Q(stg_reg[130]) );
  DFFQX1 stg_reg_reg_4__3_ ( .D(n2112), .CK(clk), .Q(stg_reg[131]) );
  DFFQX1 stg_reg_reg_4__4_ ( .D(n2111), .CK(clk), .Q(stg_reg[132]) );
  DFFX1 stg_reg_reg_1__0_ ( .D(n2243), .CK(clk), .Q(n1485), .QN(n2462) );
  DFFX1 stg_reg_reg_1__1_ ( .D(n2242), .CK(clk), .Q(n1506), .QN(n2454) );
  DFFX1 stg_reg_reg_1__2_ ( .D(n2241), .CK(clk), .Q(n1509), .QN(n2449) );
  DFFX1 stg_reg_reg_1__3_ ( .D(n2240), .CK(clk), .Q(n1512), .QN(n2444) );
  DFFX1 stg_reg_reg_1__4_ ( .D(n2239), .CK(clk), .Q(n1515), .QN(n2439) );
  DFFX1 stg_reg_reg_1__5_ ( .D(n2238), .CK(clk), .Q(n1518), .QN(n2434) );
  DFFX1 stg_reg_reg_2__0_ ( .D(n2275), .CK(clk), .Q(n1533), .QN(n3143) );
  DFFX1 stg_reg_reg_2__1_ ( .D(n2274), .CK(clk), .Q(n1554), .QN(n3138) );
  DFFX1 stg_reg_reg_2__2_ ( .D(n2273), .CK(clk), .Q(n1557), .QN(n3134) );
  DFFX1 stg_reg_reg_2__3_ ( .D(n2272), .CK(clk), .Q(n1560), .QN(n3130) );
  DFFX1 stg_reg_reg_2__4_ ( .D(n2271), .CK(clk), .Q(n1563), .QN(n3126) );
  DFFX1 stg_reg_reg_2__5_ ( .D(n2270), .CK(clk), .Q(n1566), .QN(n3121) );
  DFFX1 stg_reg_reg_0__0_ ( .D(n2211), .CK(clk), .Q(n1437), .QN(n1143) );
  DFFX1 stg_reg_reg_0__1_ ( .D(n2210), .CK(clk), .Q(n1458), .QN(n11370) );
  DFFX1 stg_reg_reg_0__2_ ( .D(n2209), .CK(clk), .Q(n1461), .QN(n11310) );
  DFFX1 stg_reg_reg_0__3_ ( .D(n2208), .CK(clk), .Q(n1464), .QN(n11250) );
  DFFX1 stg_reg_reg_0__4_ ( .D(n2207), .CK(clk), .Q(n1467), .QN(n11190) );
  DFFX1 stg_reg_reg_3__0_ ( .D(n2307), .CK(clk), .Q(n1581), .QN(n2551) );
  DFFX1 stg_reg_reg_3__1_ ( .D(n2306), .CK(clk), .Q(n1595), .QN(n2545) );
  DFFX1 stg_reg_reg_3__2_ ( .D(n2305), .CK(clk), .Q(n1597), .QN(n2539) );
  DFFX1 stg_reg_reg_3__3_ ( .D(n2304), .CK(clk), .Q(n1599), .QN(n2533) );
  DFFX1 stg_reg_reg_3__4_ ( .D(n2303), .CK(clk), .Q(n1601), .QN(n2527) );
  DFFX1 stg_reg_reg_3__5_ ( .D(n2302), .CK(clk), .Q(n1603), .QN(n2521) );
  DFFQX1 data_reg_7__0_ ( .D(data_8__0_), .CK(clk), .Q(data_7__0_) );
  DFFQX1 stg_reg_reg_15__6_ ( .D(n1870), .CK(clk), .Q(stg_reg[6]) );
  DFFQX1 stg_reg_reg_15__7_ ( .D(n1869), .CK(clk), .Q(stg_reg[7]) );
  DFFQX1 stg_reg_reg_5__0_ ( .D(n2035), .CK(clk), .Q(stg_reg[96]) );
  DFFQX1 stg_reg_reg_5__6_ ( .D(n2029), .CK(clk), .Q(stg_reg[102]) );
  DFFQX1 stg_reg_reg_5__7_ ( .D(n2028), .CK(clk), .Q(stg_reg[103]) );
  DFFQX1 stg_reg_reg_5__22_ ( .D(n2013), .CK(clk), .Q(stg_reg[118]) );
  DFFX1 stg_reg_reg_13__0_ ( .D(n2067), .CK(clk), .Q(n1487), .QN(n3061) );
  DFFX1 stg_reg_reg_9__0_ ( .D(n2099), .CK(clk), .Q(n1486), .QN(n3060) );
  DFFX1 stg_reg_reg_13__1_ ( .D(n2066), .CK(clk), .Q(n1508), .QN(n3047) );
  DFFX1 stg_reg_reg_9__1_ ( .D(n2098), .CK(clk), .Q(n1507), .QN(n3046) );
  DFFX1 stg_reg_reg_13__2_ ( .D(n2065), .CK(clk), .Q(n1511), .QN(n3034) );
  DFFX1 stg_reg_reg_9__2_ ( .D(n2097), .CK(clk), .Q(n1510), .QN(n3033) );
  DFFX1 stg_reg_reg_13__3_ ( .D(n2064), .CK(clk), .Q(n1514), .QN(n3021) );
  DFFX1 stg_reg_reg_9__3_ ( .D(n2096), .CK(clk), .Q(n1513), .QN(n3020) );
  DFFX1 stg_reg_reg_13__4_ ( .D(n2063), .CK(clk), .Q(n1517), .QN(n3008) );
  DFFX1 stg_reg_reg_9__4_ ( .D(n2095), .CK(clk), .Q(n1516), .QN(n3007) );
  DFFX1 stg_reg_reg_13__5_ ( .D(n2062), .CK(clk), .Q(n1520), .QN(n2995) );
  DFFX1 stg_reg_reg_9__5_ ( .D(n2094), .CK(clk), .Q(n1519), .QN(n2994) );
  DFFX1 stg_reg_reg_13__6_ ( .D(n2061), .CK(clk), .Q(n1523), .QN(n2982) );
  DFFX1 stg_reg_reg_9__6_ ( .D(n2093), .CK(clk), .Q(n1522), .QN(n2981) );
  DFFX1 stg_reg_reg_13__7_ ( .D(n2060), .CK(clk), .Q(n1526), .QN(n2969) );
  DFFX1 stg_reg_reg_11__16_ ( .D(n1891), .CK(clk), .Q(n1758), .QN(n2851) );
  DFFX1 stg_reg_reg_11__17_ ( .D(n1890), .CK(clk), .Q(n1772), .QN(n2841) );
  DFFX1 stg_reg_reg_11__18_ ( .D(n1889), .CK(clk), .Q(n1774), .QN(n2831) );
  DFFX1 stg_reg_reg_11__19_ ( .D(n1888), .CK(clk), .Q(n1776), .QN(n2821) );
  DFFX1 stg_reg_reg_11__20_ ( .D(n1887), .CK(clk), .Q(n1778), .QN(n2811) );
  DFFX1 stg_reg_reg_11__21_ ( .D(n1886), .CK(clk), .Q(n1780), .QN(n2801) );
  DFFX1 stg_reg_reg_11__22_ ( .D(n1885), .CK(clk), .Q(n1782), .QN(n2791) );
  DFFX1 stg_reg_reg_11__23_ ( .D(n1884), .CK(clk), .Q(n1784), .QN(n2781) );
  DFFX1 stg_reg_reg_14__16_ ( .D(n1955), .CK(clk), .Q(n1711), .QN(n2852) );
  DFFX1 stg_reg_reg_14__17_ ( .D(n1954), .CK(clk), .Q(n1732), .QN(n2842) );
  DFFX1 stg_reg_reg_14__18_ ( .D(n1953), .CK(clk), .Q(n1735), .QN(n2832) );
  DFFX1 stg_reg_reg_14__19_ ( .D(n1952), .CK(clk), .Q(n1738), .QN(n2822) );
  DFFX1 stg_reg_reg_14__20_ ( .D(n1951), .CK(clk), .Q(n1741), .QN(n2812) );
  DFFX1 stg_reg_reg_14__21_ ( .D(n1950), .CK(clk), .Q(n1744), .QN(n2802) );
  DFFX1 stg_reg_reg_14__22_ ( .D(n1949), .CK(clk), .Q(n1747), .QN(n2792) );
  DFFX1 stg_reg_reg_13__16_ ( .D(n2051), .CK(clk), .Q(n1663), .QN(n2854) );
  DFFX1 stg_reg_reg_9__16_ ( .D(n2083), .CK(clk), .Q(n1662), .QN(n2853) );
  DFFX1 stg_reg_reg_13__17_ ( .D(n2050), .CK(clk), .Q(n1684), .QN(n2844) );
  DFFX1 stg_reg_reg_9__17_ ( .D(n2082), .CK(clk), .Q(n1683), .QN(n2843) );
  DFFX1 stg_reg_reg_13__18_ ( .D(n2049), .CK(clk), .Q(n1687), .QN(n2834) );
  DFFX1 stg_reg_reg_9__18_ ( .D(n2081), .CK(clk), .Q(n1686), .QN(n2833) );
  DFFX1 stg_reg_reg_13__19_ ( .D(n2048), .CK(clk), .Q(n1690), .QN(n2824) );
  DFFX1 stg_reg_reg_9__19_ ( .D(n2080), .CK(clk), .Q(n1689), .QN(n2823) );
  DFFX1 stg_reg_reg_13__20_ ( .D(n2047), .CK(clk), .Q(n1693), .QN(n2814) );
  DFFX1 stg_reg_reg_9__20_ ( .D(n2079), .CK(clk), .Q(n1692), .QN(n2813) );
  DFFX1 stg_reg_reg_13__21_ ( .D(n2046), .CK(clk), .Q(n1696), .QN(n2804) );
  DFFX1 stg_reg_reg_9__21_ ( .D(n2078), .CK(clk), .Q(n1695), .QN(n2803) );
  DFFX1 stg_reg_reg_13__22_ ( .D(n2045), .CK(clk), .Q(n1699), .QN(n2794) );
  DFFX1 stg_reg_reg_9__22_ ( .D(n2077), .CK(clk), .Q(n1698), .QN(n2793) );
  DFFX1 stg_reg_reg_9__23_ ( .D(n2076), .CK(clk), .Q(n1701), .QN(n2783) );
  DFFX1 stg_reg_reg_14__0_ ( .D(n1971), .CK(clk), .Q(n1535), .QN(n3147) );
  DFFX1 stg_reg_reg_14__1_ ( .D(n1970), .CK(clk), .Q(n1556), .QN(n3141) );
  DFFX1 stg_reg_reg_14__2_ ( .D(n1969), .CK(clk), .Q(n1559), .QN(n3137) );
  DFFX1 stg_reg_reg_14__3_ ( .D(n1968), .CK(clk), .Q(n1562), .QN(n3133) );
  DFFX1 stg_reg_reg_14__4_ ( .D(n1967), .CK(clk), .Q(n1565), .QN(n3129) );
  DFFX1 stg_reg_reg_14__5_ ( .D(n1966), .CK(clk), .Q(n1568), .QN(n3125) );
  DFFX1 stg_reg_reg_14__6_ ( .D(n1965), .CK(clk), .Q(n1571), .QN(n3120) );
  DFFX1 stg_reg_reg_14__7_ ( .D(n1964), .CK(clk), .Q(n1574), .QN(n3115) );
  DFFX1 stg_reg_reg_11__0_ ( .D(n1907), .CK(clk), .Q(n1582), .QN(n3059) );
  DFFX1 stg_reg_reg_11__1_ ( .D(n1906), .CK(clk), .Q(n1596), .QN(n3045) );
  DFFX1 stg_reg_reg_11__2_ ( .D(n1905), .CK(clk), .Q(n1598), .QN(n3032) );
  DFFX1 stg_reg_reg_11__3_ ( .D(n1904), .CK(clk), .Q(n1600), .QN(n3019) );
  DFFX1 stg_reg_reg_11__4_ ( .D(n1903), .CK(clk), .Q(n1602), .QN(n3006) );
  DFFX1 stg_reg_reg_11__5_ ( .D(n1902), .CK(clk), .Q(n1604), .QN(n2993) );
  DFFX1 stg_reg_reg_11__6_ ( .D(n1901), .CK(clk), .Q(n1606), .QN(n2980) );
  DFFQX1 stg_reg_reg_6__16_ ( .D(n1923), .CK(clk), .Q(stg_reg[80]) );
  DFFQX1 stg_reg_reg_6__18_ ( .D(n1921), .CK(clk), .Q(stg_reg[82]) );
  DFFQX1 stg_reg_reg_6__20_ ( .D(n1919), .CK(clk), .Q(stg_reg[84]) );
  DFFQX1 stg_reg_reg_6__23_ ( .D(n1916), .CK(clk), .Q(stg_reg[87]) );
  DFFQX1 stg_reg_reg_7__16_ ( .D(n1828), .CK(clk), .Q(stg_reg[48]) );
  DFFQX1 stg_reg_reg_7__18_ ( .D(n1826), .CK(clk), .Q(stg_reg[50]) );
  DFFQX1 stg_reg_reg_7__20_ ( .D(n1824), .CK(clk), .Q(stg_reg[52]) );
  DFFQX1 stg_reg_reg_7__21_ ( .D(n1823), .CK(clk), .Q(stg_reg[53]) );
  DFFQX1 stg_reg_reg_7__0_ ( .D(n1844), .CK(clk), .Q(stg_reg[32]) );
  DFFQX1 stg_reg_reg_7__2_ ( .D(n1842), .CK(clk), .Q(stg_reg[34]) );
  DFFQX1 stg_reg_reg_7__4_ ( .D(n1840), .CK(clk), .Q(stg_reg[36]) );
  DFFQX1 stg_reg_reg_7__5_ ( .D(n1839), .CK(clk), .Q(stg_reg[37]) );
  DFFQX1 stg_reg_reg_6__0_ ( .D(n1939), .CK(clk), .Q(stg_reg[64]) );
  DFFQX1 stg_reg_reg_6__2_ ( .D(n1937), .CK(clk), .Q(stg_reg[66]) );
  DFFQX1 stg_reg_reg_6__4_ ( .D(n1935), .CK(clk), .Q(stg_reg[68]) );
  DFFQX1 stg_reg_reg_6__6_ ( .D(n1933), .CK(clk), .Q(stg_reg[70]) );
  DFFQX1 stg_reg_reg_6__7_ ( .D(n1932), .CK(clk), .Q(stg_reg[71]) );
  DFFX1 stg_reg_reg_10__16_ ( .D(n1987), .CK(clk), .Q(n1710), .QN(n98) );
  DFFX1 stg_reg_reg_10__17_ ( .D(n1986), .CK(clk), .Q(n1731), .QN(n116) );
  DFFX1 stg_reg_reg_10__18_ ( .D(n1985), .CK(clk), .Q(n1734), .QN(n115) );
  DFFX1 stg_reg_reg_10__19_ ( .D(n1984), .CK(clk), .Q(n1737), .QN(n119) );
  DFFX1 stg_reg_reg_10__20_ ( .D(n1983), .CK(clk), .Q(n1740), .QN(n118) );
  DFFX1 stg_reg_reg_10__21_ ( .D(n1982), .CK(clk), .Q(n1743), .QN(n117) );
  DFFX1 stg_reg_reg_10__23_ ( .D(n1980), .CK(clk), .Q(n1749), .QN(n125) );
  DFFX1 stg_reg_reg_10__0_ ( .D(n2003), .CK(clk), .Q(n1534), .QN(n114) );
  DFFX1 stg_reg_reg_10__1_ ( .D(n2002), .CK(clk), .Q(n1555), .QN(n100) );
  DFFX1 stg_reg_reg_10__2_ ( .D(n2001), .CK(clk), .Q(n1558), .QN(n99) );
  DFFX1 stg_reg_reg_10__3_ ( .D(n2000), .CK(clk), .Q(n1561), .QN(n102) );
  DFFX1 stg_reg_reg_10__4_ ( .D(n1999), .CK(clk), .Q(n1564), .QN(n101) );
  DFFX1 stg_reg_reg_10__5_ ( .D(n1998), .CK(clk), .Q(n1567), .QN(n3124) );
  DFFRX2 cnt_reg_3_ ( .D(N38), .CK(clk), .RN(n3149), .Q(mul_2_Wn[13]), .QN(
        n1810) );
  DFFQX1 data_reg_12__0_ ( .D(data_13__0_), .CK(clk), .Q(data_12__0_) );
  DFFQX1 data_reg_1__0_ ( .D(data_2__0_), .CK(clk), .Q(data_1__0_) );
  DFFQX1 data_reg_14__0_ ( .D(fir_d[0]), .CK(clk), .Q(data_14__0_) );
  DFFQX1 data_reg_13__0_ ( .D(data_14__0_), .CK(clk), .Q(data_13__0_) );
  DFFQX1 data_reg_3__0_ ( .D(data_4__0_), .CK(clk), .Q(data_3__0_) );
  DFFQX1 data_reg_2__0_ ( .D(data_3__0_), .CK(clk), .Q(data_2__0_) );
  DFFXL stg_reg_reg_9__13_ ( .D(n2086), .CK(clk), .Q(n1498), .QN(n93) );
  DFFQXL stg_reg_reg_15__13_ ( .D(n1863), .CK(clk), .Q(stg_reg[13]) );
  DFFQXL stg_reg_reg_15__28_ ( .D(n1848), .CK(clk), .Q(stg_reg[28]) );
  DFFQXL stg_reg_reg_15__27_ ( .D(n1849), .CK(clk), .Q(stg_reg[27]) );
  DFFQXL stg_reg_reg_15__12_ ( .D(n1864), .CK(clk), .Q(stg_reg[12]) );
  DFFQXL stg_reg_reg_15__11_ ( .D(n1865), .CK(clk), .Q(stg_reg[11]) );
  DFFQXL stg_reg_reg_15__26_ ( .D(n1850), .CK(clk), .Q(stg_reg[26]) );
  DFFQXL stg_reg_reg_15__10_ ( .D(n1866), .CK(clk), .Q(stg_reg[10]) );
  DFFQXL stg_reg_reg_15__22_ ( .D(n1854), .CK(clk), .Q(stg_reg[22]) );
  DFFQXL stg_reg_reg_15__24_ ( .D(n1852), .CK(clk), .Q(stg_reg[24]) );
  DFFQXL stg_reg_reg_15__8_ ( .D(n1868), .CK(clk), .Q(stg_reg[8]) );
  DFFQXL stg_reg_reg_15__25_ ( .D(n1851), .CK(clk), .Q(stg_reg[25]) );
  DFFQXL stg_reg_reg_15__9_ ( .D(n1867), .CK(clk), .Q(stg_reg[9]) );
  DFFQXL stg_reg_reg_15__23_ ( .D(n1853), .CK(clk), .Q(stg_reg[23]) );
  DFFQXL stg_reg_reg_5__27_ ( .D(n2008), .CK(clk), .Q(stg_reg[123]) );
  DFFQXL stg_reg_reg_5__28_ ( .D(n2007), .CK(clk), .Q(stg_reg[124]) );
  DFFQXL stg_reg_reg_5__11_ ( .D(n2024), .CK(clk), .Q(stg_reg[107]) );
  DFFQXL stg_reg_reg_5__12_ ( .D(n2023), .CK(clk), .Q(stg_reg[108]) );
  DFFQXL stg_reg_reg_5__26_ ( .D(n2009), .CK(clk), .Q(stg_reg[122]) );
  DFFQXL stg_reg_reg_5__10_ ( .D(n2025), .CK(clk), .Q(stg_reg[106]) );
  DFFQXL stg_reg_reg_5__24_ ( .D(n2011), .CK(clk), .Q(stg_reg[120]) );
  DFFQXL stg_reg_reg_5__8_ ( .D(n2027), .CK(clk), .Q(stg_reg[104]) );
  DFFQXL stg_reg_reg_5__25_ ( .D(n2010), .CK(clk), .Q(stg_reg[121]) );
  DFFQXL stg_reg_reg_5__9_ ( .D(n2026), .CK(clk), .Q(stg_reg[105]) );
  DFFQXL stg_reg_reg_7__8_ ( .D(n1836), .CK(clk), .Q(stg_reg[40]) );
  DFFQXL stg_reg_reg_6__8_ ( .D(n1931), .CK(clk), .Q(stg_reg[72]) );
  DFFRX4 cnt_reg_2_ ( .D(N37), .CK(clk), .RN(n3149), .Q(n176), .QN(n1790) );
  DFFRX4 cnt_reg_0_ ( .D(n842), .CK(clk), .RN(n3149), .Q(n177), .QN(n1789) );
  DFFX1 stg_reg_reg_10__22_ ( .D(n1981), .CK(clk), .Q(n1746), .QN(n126) );
  DFFQX1 stg_reg_reg_7__22_ ( .D(n1822), .CK(clk), .Q(stg_reg[54]) );
  DFFQX1 stg_reg_reg_7__23_ ( .D(n1821), .CK(clk), .Q(stg_reg[55]) );
  DFFQX1 stg_reg_reg_7__6_ ( .D(n1838), .CK(clk), .Q(stg_reg[38]) );
  DFFQX1 stg_reg_reg_7__7_ ( .D(n1837), .CK(clk), .Q(stg_reg[39]) );
  DFFQX1 stg_reg_reg_6__22_ ( .D(n1917), .CK(clk), .Q(stg_reg[86]) );
  DFFQX1 stg_reg_reg_15__16_ ( .D(n1860), .CK(clk), .Q(stg_reg[16]) );
  DFFXL stg_reg_reg_13__14_ ( .D(n2053), .CK(clk), .Q(n1502), .QN(n110) );
  DFFXL stg_reg_reg_9__14_ ( .D(n2085), .CK(clk), .Q(n1501), .QN(n95) );
  DFFXL stg_reg_reg_9__15_ ( .D(n2084), .CK(clk), .Q(n1504) );
  DFFXL stg_reg_reg_9__30_ ( .D(n2069), .CK(clk), .Q(n1677), .QN(n92) );
  DFFXL stg_reg_reg_11__31_ ( .D(n1876), .CK(clk), .Q(n1770), .QN(n90) );
  DFFXL stg_reg_reg_14__31_ ( .D(n1940), .CK(clk), .Q(n1729), .QN(n89) );
  DFFXL stg_reg_reg_13__31_ ( .D(n2036), .CK(clk), .Q(n1681), .QN(n91) );
  DFFXL stg_reg_reg_9__31_ ( .D(n2068), .CK(clk), .Q(n1680), .QN(n96) );
  DFFXL stg_reg_reg_14__14_ ( .D(n1957), .CK(clk), .Q(n1550), .QN(n94) );
  DFFXL stg_reg_reg_11__13_ ( .D(n1894), .CK(clk), .Q(n1590), .QN(n108) );
  DFFXL stg_reg_reg_11__14_ ( .D(n1893), .CK(clk), .Q(n1592), .QN(n112) );
  DFFXL stg_reg_reg_11__15_ ( .D(n1892), .CK(clk), .Q(n1594), .QN(n111) );
  DFFXL stg_reg_reg_13__15_ ( .D(n2052), .CK(clk), .Q(n1505), .QN(n113) );
  DFFXL stg_reg_reg_14__15_ ( .D(n1956), .CK(clk), .Q(n1553), .QN(n97) );
  DFFQXL stg_reg_reg_15__30_ ( .D(n1846), .CK(clk), .Q(stg_reg[30]) );
  DFFQXL stg_reg_reg_15__14_ ( .D(n1862), .CK(clk), .Q(stg_reg[14]) );
  DFFQXL stg_reg_reg_15__31_ ( .D(n1845), .CK(clk), .Q(stg_reg[31]) );
  DFFQXL stg_reg_reg_15__15_ ( .D(n1861), .CK(clk), .Q(stg_reg[15]) );
  DFFQXL stg_reg_reg_5__13_ ( .D(n2022), .CK(clk), .Q(stg_reg[109]) );
  DFFQXL stg_reg_reg_5__14_ ( .D(n2021), .CK(clk), .Q(stg_reg[110]) );
  DFFQXL stg_reg_reg_5__29_ ( .D(n2006), .CK(clk), .Q(stg_reg[125]) );
  DFFQXL stg_reg_reg_5__30_ ( .D(n2005), .CK(clk), .Q(stg_reg[126]) );
  DFFQXL stg_reg_reg_5__15_ ( .D(n2020), .CK(clk), .Q(stg_reg[111]) );
  DFFQXL stg_reg_reg_5__31_ ( .D(n2004), .CK(clk), .Q(stg_reg[127]) );
  DFFXL stg_reg_reg_10__31_ ( .D(n1972), .CK(clk), .Q(n1728), .QN(n152) );
  DFFXL stg_reg_reg_10__15_ ( .D(n1988), .CK(clk), .Q(n1552), .QN(n150) );
  DFFQXL stg_reg_reg_7__11_ ( .D(n1833), .CK(clk), .Q(stg_reg[43]) );
  DFFQXL stg_reg_reg_7__26_ ( .D(n1818), .CK(clk), .Q(stg_reg[58]) );
  DFFQXL stg_reg_reg_7__10_ ( .D(n1834), .CK(clk), .Q(stg_reg[42]) );
  DFFQXL stg_reg_reg_6__10_ ( .D(n1929), .CK(clk), .Q(stg_reg[74]) );
  DFFQXL stg_reg_reg_6__28_ ( .D(n1911), .CK(clk), .Q(stg_reg[92]) );
  DFFQXL stg_reg_reg_6__26_ ( .D(n1913), .CK(clk), .Q(stg_reg[90]) );
  DFFQXL stg_reg_reg_7__28_ ( .D(n1816), .CK(clk), .Q(stg_reg[60]) );
  DFFQXL stg_reg_reg_7__30_ ( .D(n1814), .CK(clk), .Q(stg_reg[62]) );
  DFFQXL stg_reg_reg_7__14_ ( .D(n1830), .CK(clk), .Q(stg_reg[46]) );
  DFFQXL stg_reg_reg_7__15_ ( .D(n1829), .CK(clk), .Q(stg_reg[47]) );
  DFFQXL stg_reg_reg_7__31_ ( .D(n1813), .CK(clk), .Q(stg_reg[63]) );
  DFFQXL stg_reg_reg_6__15_ ( .D(n1924), .CK(clk), .Q(stg_reg[79]) );
  DFFQXL stg_reg_reg_6__30_ ( .D(n1909), .CK(clk), .Q(stg_reg[94]) );
  DFFQXL stg_reg_reg_6__31_ ( .D(n1908), .CK(clk), .Q(stg_reg[95]) );
  DFFX1 stg_reg_reg_10__24_ ( .D(n1979), .CK(clk), .Q(n1752), .QN(n124) );
  DFFXL stg_reg_reg_10__13_ ( .D(n1990), .CK(clk), .Q(n1546), .QN(n132) );
  DFFXL stg_reg_reg_10__14_ ( .D(n1989), .CK(clk), .Q(n1549), .QN(n151) );
  DFFQXL stg_reg_reg_6__13_ ( .D(n1926), .CK(clk), .Q(stg_reg[77]) );
  DFFQXL stg_reg_reg_6__12_ ( .D(n1927), .CK(clk), .Q(stg_reg[76]) );
  DFFQXL stg_reg_reg_7__27_ ( .D(n1817), .CK(clk), .Q(stg_reg[59]) );
  DFFQXL stg_reg_reg_7__29_ ( .D(n1815), .CK(clk), .Q(stg_reg[61]) );
  DFFQXL stg_reg_reg_7__12_ ( .D(n1832), .CK(clk), .Q(stg_reg[44]) );
  DFFQXL stg_reg_reg_7__13_ ( .D(n1831), .CK(clk), .Q(stg_reg[45]) );
  DFFQXL stg_reg_reg_6__14_ ( .D(n1925), .CK(clk), .Q(stg_reg[78]) );
  DFFQX1 stg_reg_reg_5__16_ ( .D(n2019), .CK(clk), .Q(stg_reg[112]) );
  DFFQX1 stg_reg_reg_15__19_ ( .D(n1857), .CK(clk), .Q(stg_reg[19]) );
  DFFQX1 stg_reg_reg_15__21_ ( .D(n1855), .CK(clk), .Q(stg_reg[21]) );
  DFFQX1 stg_reg_reg_15__5_ ( .D(n1871), .CK(clk), .Q(stg_reg[5]) );
  DFFQX1 stg_reg_reg_5__21_ ( .D(n2014), .CK(clk), .Q(stg_reg[117]) );
  DFFQXL stg_reg_reg_7__24_ ( .D(n1820), .CK(clk), .Q(stg_reg[56]) );
  DFFQXL stg_reg_reg_6__11_ ( .D(n1928), .CK(clk), .Q(stg_reg[75]) );
  DFFQXL stg_reg_reg_6__29_ ( .D(n1910), .CK(clk), .Q(stg_reg[93]) );
  DFFQXL stg_reg_reg_6__27_ ( .D(n1912), .CK(clk), .Q(stg_reg[91]) );
  DFFQX1 stg_reg_reg_5__5_ ( .D(n2030), .CK(clk), .Q(stg_reg[101]) );
  DFFQX1 stg_reg_reg_5__20_ ( .D(n2015), .CK(clk), .Q(stg_reg[116]) );
  DFFQX1 stg_reg_reg_6__21_ ( .D(n1918), .CK(clk), .Q(stg_reg[85]) );
  DFFQXL stg_reg_reg_7__9_ ( .D(n1835), .CK(clk), .Q(stg_reg[41]) );
  DFFQXL stg_reg_reg_6__9_ ( .D(n1930), .CK(clk), .Q(stg_reg[73]) );
  DFFQX1 stg_reg_reg_15__20_ ( .D(n1856), .CK(clk), .Q(stg_reg[20]) );
  DFFQX1 stg_reg_reg_15__4_ ( .D(n1872), .CK(clk), .Q(stg_reg[4]) );
  DFFQX1 stg_reg_reg_5__4_ ( .D(n2031), .CK(clk), .Q(stg_reg[100]) );
  DFFX1 stg_reg_reg_10__7_ ( .D(n1996), .CK(clk), .Q(n1573), .QN(n105) );
  DFFQX1 stg_reg_reg_6__5_ ( .D(n1934), .CK(clk), .Q(stg_reg[69]) );
  DFFQX1 fft_d0_reg_15_ ( .D(N678), .CK(clk), .Q(n3719) );
  DFFQX1 fft_d0_reg_31_ ( .D(N694), .CK(clk), .Q(n3707) );
  DFFRX1 fft_valid_reg ( .D(N39), .CK(clk), .RN(n3149), .QN(n7160) );
  MDFFHQX1 fft_d2_reg_0_ ( .D0(stg_reg[128]), .D1(fft_d3[0]), .S0(n10240), 
        .CK(clk), .Q(n3290) );
  MDFFHQX1 fft_d10_reg_0_ ( .D0(stg_reg[96]), .D1(fft_d11[0]), .S0(n10330), 
        .CK(clk), .Q(n3546) );
  MDFFHQX1 fft_d10_reg_2_ ( .D0(stg_reg[98]), .D1(fft_d11[2]), .S0(n10320), 
        .CK(clk), .Q(n3544) );
  DFFQX1 stg_reg_reg_5__2_ ( .D(n2033), .CK(clk), .Q(stg_reg[98]) );
  MDFFHQX1 fft_d10_reg_4_ ( .D0(stg_reg[100]), .D1(fft_d11[4]), .S0(n10310), 
        .CK(clk), .Q(n3542) );
  MDFFHQX1 fft_d10_reg_6_ ( .D0(stg_reg[102]), .D1(fft_d11[6]), .S0(n10300), 
        .CK(clk), .Q(n3540) );
  MDFFHQX1 fft_d10_reg_8_ ( .D0(stg_reg[104]), .D1(fft_d11[8]), .S0(n10290), 
        .CK(clk), .Q(n3538) );
  MDFFHQX1 fft_d10_reg_10_ ( .D0(stg_reg[106]), .D1(fft_d11[10]), .S0(n10280), 
        .CK(clk), .Q(n3536) );
  MDFFHQX1 fft_d10_reg_12_ ( .D0(stg_reg[108]), .D1(fft_d11[12]), .S0(n10270), 
        .CK(clk), .Q(n3534) );
  MDFFHQX1 fft_d10_reg_14_ ( .D0(stg_reg[110]), .D1(fft_d11[14]), .S0(n10260), 
        .CK(clk), .Q(n3532) );
  MDFFHQX1 fft_d6_reg_16_ ( .D0(stg_reg[80]), .D1(fft_d7[16]), .S0(n10250), 
        .CK(clk), .Q(n3402) );
  MDFFHQX1 fft_d6_reg_18_ ( .D0(stg_reg[82]), .D1(fft_d7[18]), .S0(n10240), 
        .CK(clk), .Q(n3400) );
  MDFFHQX1 fft_d6_reg_20_ ( .D0(stg_reg[84]), .D1(fft_d7[20]), .S0(n10230), 
        .CK(clk), .Q(n3398) );
  MDFFHQX1 fft_d6_reg_22_ ( .D0(stg_reg[86]), .D1(fft_d7[22]), .S0(n10220), 
        .CK(clk), .Q(n3396) );
  MDFFHQX1 fft_d6_reg_24_ ( .D0(stg_reg[88]), .D1(fft_d7[24]), .S0(n10210), 
        .CK(clk), .Q(n3394) );
  DFFQXL stg_reg_reg_6__24_ ( .D(n1915), .CK(clk), .Q(stg_reg[88]) );
  MDFFHQX1 fft_d6_reg_26_ ( .D0(stg_reg[90]), .D1(fft_d7[26]), .S0(n10200), 
        .CK(clk), .Q(n3392) );
  MDFFHQX1 fft_d6_reg_28_ ( .D0(stg_reg[92]), .D1(fft_d7[28]), .S0(n10190), 
        .CK(clk), .Q(n3390) );
  MDFFHQX1 fft_d10_reg_29_ ( .D0(stg_reg[125]), .D1(fft_d11[29]), .S0(n10180), 
        .CK(clk), .Q(n3517) );
  MDFFHQX1 fft_d14_reg_29_ ( .D0(stg_reg[61]), .D1(fft_d15[29]), .S0(n10170), 
        .CK(clk), .Q(n3645) );
  MDFFHQX1 fft_d2_reg_30_ ( .D0(stg_reg[158]), .D1(fft_d3[30]), .S0(n10160), 
        .CK(clk), .Q(n3260) );
  MDFFHQX1 fft_d6_reg_30_ ( .D0(stg_reg[94]), .D1(fft_d7[30]), .S0(n10150), 
        .CK(clk), .Q(n3388) );
  MDFFHQX1 fft_d10_reg_30_ ( .D0(stg_reg[126]), .D1(fft_d11[30]), .S0(n10140), 
        .CK(clk), .Q(n3516) );
  MDFFHQX1 fft_d14_reg_30_ ( .D0(stg_reg[62]), .D1(fft_d15[30]), .S0(n10130), 
        .CK(clk), .Q(n3644) );
  MDFFHQX1 fft_d2_reg_31_ ( .D0(stg_reg[159]), .D1(fft_d3[31]), .S0(n10120), 
        .CK(clk), .Q(n3259) );
  MDFFHQX1 fft_d6_reg_31_ ( .D0(stg_reg[95]), .D1(fft_d7[31]), .S0(n10110), 
        .CK(clk), .Q(n3387) );
  MDFFHQX1 fft_d10_reg_31_ ( .D0(stg_reg[127]), .D1(fft_d11[31]), .S0(n10240), 
        .CK(clk), .Q(n3515) );
  DFFQX1 fft_d7_reg_0_ ( .D(N1111), .CK(clk), .Q(n3450) );
  DFFQX1 fft_d15_reg_0_ ( .D(stg_reg[0]), .CK(clk), .Q(n3706) );
  DFFQX1 fft_d3_reg_1_ ( .D(N1048), .CK(clk), .Q(n3321) );
  DFFQX1 fft_d7_reg_1_ ( .D(N1112), .CK(clk), .Q(n3449) );
  DFFQX1 fft_d11_reg_1_ ( .D(N1080), .CK(clk), .Q(n3577) );
  DFFQX1 fft_d15_reg_1_ ( .D(stg_reg[1]), .CK(clk), .Q(n3705) );
  DFFQX1 fft_d3_reg_2_ ( .D(N1049), .CK(clk), .Q(n3320) );
  DFFQX1 fft_d7_reg_2_ ( .D(N1113), .CK(clk), .Q(n3448) );
  DFFQX1 fft_d15_reg_2_ ( .D(stg_reg[2]), .CK(clk), .Q(n3704) );
  DFFQX1 fft_d3_reg_3_ ( .D(N1050), .CK(clk), .Q(n3319) );
  DFFQX1 fft_d7_reg_3_ ( .D(N1114), .CK(clk), .Q(n3447) );
  DFFQX1 fft_d11_reg_3_ ( .D(N1082), .CK(clk), .Q(n3575) );
  DFFQX1 fft_d15_reg_3_ ( .D(stg_reg[3]), .CK(clk), .Q(n3703) );
  DFFQX1 fft_d3_reg_4_ ( .D(N1051), .CK(clk), .Q(n3318) );
  DFFQX1 fft_d7_reg_4_ ( .D(N1115), .CK(clk), .Q(n3446) );
  DFFQX1 fft_d15_reg_4_ ( .D(stg_reg[4]), .CK(clk), .Q(n3702) );
  DFFQX1 fft_d3_reg_5_ ( .D(N1052), .CK(clk), .Q(n3317) );
  DFFQX1 fft_d7_reg_5_ ( .D(N1116), .CK(clk), .Q(n3445) );
  DFFQX1 fft_d11_reg_5_ ( .D(N1084), .CK(clk), .Q(n3573) );
  DFFQX1 fft_d15_reg_5_ ( .D(stg_reg[5]), .CK(clk), .Q(n3701) );
  DFFQX1 fft_d3_reg_6_ ( .D(N1053), .CK(clk), .Q(n3316) );
  DFFQX1 fft_d7_reg_6_ ( .D(N1117), .CK(clk), .Q(n3444) );
  DFFQX1 fft_d15_reg_6_ ( .D(stg_reg[6]), .CK(clk), .Q(n3700) );
  DFFQX1 fft_d3_reg_7_ ( .D(N1054), .CK(clk), .Q(n3315) );
  DFFQX1 fft_d7_reg_7_ ( .D(N1118), .CK(clk), .Q(n3443) );
  DFFQX1 fft_d11_reg_7_ ( .D(N1086), .CK(clk), .Q(n3571) );
  DFFQX1 fft_d15_reg_7_ ( .D(stg_reg[7]), .CK(clk), .Q(n3699) );
  DFFQX1 fft_d3_reg_8_ ( .D(N1055), .CK(clk), .Q(n3314) );
  DFFQX1 fft_d7_reg_8_ ( .D(N1119), .CK(clk), .Q(n3442) );
  DFFQX1 fft_d15_reg_8_ ( .D(stg_reg[8]), .CK(clk), .Q(n3698) );
  DFFQX1 fft_d3_reg_9_ ( .D(N1056), .CK(clk), .Q(n3313) );
  DFFQX1 fft_d7_reg_9_ ( .D(N1120), .CK(clk), .Q(n3441) );
  DFFQX1 fft_d11_reg_9_ ( .D(N1088), .CK(clk), .Q(n3569) );
  DFFQX1 fft_d15_reg_9_ ( .D(stg_reg[9]), .CK(clk), .Q(n3697) );
  DFFQX1 fft_d3_reg_10_ ( .D(N1057), .CK(clk), .Q(n3312) );
  DFFQX1 fft_d7_reg_10_ ( .D(N1121), .CK(clk), .Q(n3440) );
  DFFQX1 fft_d15_reg_10_ ( .D(stg_reg[10]), .CK(clk), .Q(n3696) );
  DFFQX1 fft_d3_reg_11_ ( .D(N1058), .CK(clk), .Q(n3311) );
  DFFQX1 fft_d7_reg_11_ ( .D(N1122), .CK(clk), .Q(n3439) );
  DFFQX1 fft_d11_reg_11_ ( .D(N1090), .CK(clk), .Q(n3567) );
  DFFQX1 fft_d15_reg_11_ ( .D(stg_reg[11]), .CK(clk), .Q(n3695) );
  DFFQX1 fft_d3_reg_12_ ( .D(N1059), .CK(clk), .Q(n3310) );
  DFFQX1 fft_d7_reg_12_ ( .D(N1123), .CK(clk), .Q(n3438) );
  DFFQX1 fft_d15_reg_12_ ( .D(stg_reg[12]), .CK(clk), .Q(n3694) );
  DFFQX1 fft_d3_reg_13_ ( .D(N1060), .CK(clk), .Q(n3309) );
  DFFQX1 fft_d7_reg_13_ ( .D(N1124), .CK(clk), .Q(n3437) );
  DFFQX1 fft_d11_reg_13_ ( .D(N1092), .CK(clk), .Q(n3565) );
  DFFQX1 fft_d15_reg_13_ ( .D(stg_reg[13]), .CK(clk), .Q(n3693) );
  DFFQX1 fft_d3_reg_14_ ( .D(N1061), .CK(clk), .Q(n3308) );
  DFFQX1 fft_d7_reg_14_ ( .D(N1125), .CK(clk), .Q(n3436) );
  DFFQX1 fft_d15_reg_14_ ( .D(stg_reg[14]), .CK(clk), .Q(n3692) );
  DFFQX1 fft_d3_reg_15_ ( .D(N1062), .CK(clk), .Q(n3307) );
  DFFQX1 fft_d7_reg_15_ ( .D(N1126), .CK(clk), .Q(n3435) );
  DFFQX1 fft_d11_reg_15_ ( .D(N1094), .CK(clk), .Q(n3563) );
  DFFQX1 fft_d15_reg_15_ ( .D(stg_reg[15]), .CK(clk), .Q(n3691) );
  DFFQX1 fft_d3_reg_16_ ( .D(N1063), .CK(clk), .Q(n3306) );
  DFFQX1 fft_d11_reg_16_ ( .D(N1095), .CK(clk), .Q(n3562) );
  DFFQX1 fft_d15_reg_16_ ( .D(stg_reg[16]), .CK(clk), .Q(n3690) );
  DFFQX1 fft_d3_reg_17_ ( .D(N1064), .CK(clk), .Q(n3305) );
  DFFQX1 fft_d7_reg_17_ ( .D(N1128), .CK(clk), .Q(n3433) );
  DFFQX1 fft_d11_reg_17_ ( .D(N1096), .CK(clk), .Q(n3561) );
  DFFQX1 fft_d15_reg_17_ ( .D(stg_reg[17]), .CK(clk), .Q(n3689) );
  DFFQX1 fft_d3_reg_18_ ( .D(N1065), .CK(clk), .Q(n3304) );
  DFFQX1 fft_d11_reg_18_ ( .D(N1097), .CK(clk), .Q(n3560) );
  DFFQX1 fft_d15_reg_18_ ( .D(stg_reg[18]), .CK(clk), .Q(n3688) );
  DFFQX1 fft_d3_reg_19_ ( .D(N1066), .CK(clk), .Q(n3303) );
  DFFQX1 fft_d7_reg_19_ ( .D(N1130), .CK(clk), .Q(n3431) );
  DFFQX1 fft_d11_reg_19_ ( .D(N1098), .CK(clk), .Q(n3559) );
  DFFQX1 fft_d15_reg_19_ ( .D(stg_reg[19]), .CK(clk), .Q(n3687) );
  DFFQX1 fft_d3_reg_20_ ( .D(N1067), .CK(clk), .Q(n3302) );
  DFFQX1 fft_d11_reg_20_ ( .D(N1099), .CK(clk), .Q(n3558) );
  DFFQX1 fft_d15_reg_20_ ( .D(stg_reg[20]), .CK(clk), .Q(n3686) );
  DFFQX1 fft_d3_reg_21_ ( .D(N1068), .CK(clk), .Q(n3301) );
  DFFQX1 fft_d7_reg_21_ ( .D(N1132), .CK(clk), .Q(n3429) );
  DFFQX1 fft_d11_reg_21_ ( .D(N1100), .CK(clk), .Q(n3557) );
  DFFQX1 fft_d15_reg_21_ ( .D(stg_reg[21]), .CK(clk), .Q(n3685) );
  DFFQX1 fft_d3_reg_22_ ( .D(N1069), .CK(clk), .Q(n3300) );
  DFFQX1 fft_d11_reg_22_ ( .D(N1101), .CK(clk), .Q(n3556) );
  DFFQX1 fft_d15_reg_22_ ( .D(stg_reg[22]), .CK(clk), .Q(n3684) );
  DFFQX1 fft_d3_reg_23_ ( .D(N1070), .CK(clk), .Q(n3299) );
  DFFQX1 fft_d7_reg_23_ ( .D(N1134), .CK(clk), .Q(n3427) );
  DFFQX1 fft_d11_reg_23_ ( .D(N1102), .CK(clk), .Q(n3555) );
  DFFQX1 fft_d15_reg_23_ ( .D(stg_reg[23]), .CK(clk), .Q(n3683) );
  DFFQX1 fft_d3_reg_24_ ( .D(N1071), .CK(clk), .Q(n3298) );
  DFFQX1 fft_d11_reg_24_ ( .D(N1103), .CK(clk), .Q(n3554) );
  DFFQX1 fft_d15_reg_24_ ( .D(stg_reg[24]), .CK(clk), .Q(n3682) );
  DFFQX1 fft_d3_reg_25_ ( .D(N1072), .CK(clk), .Q(n3297) );
  DFFQX1 fft_d7_reg_25_ ( .D(N1136), .CK(clk), .Q(n3425) );
  DFFQX1 fft_d11_reg_25_ ( .D(N1104), .CK(clk), .Q(n3553) );
  DFFQX1 fft_d15_reg_25_ ( .D(stg_reg[25]), .CK(clk), .Q(n3681) );
  DFFQX1 fft_d3_reg_26_ ( .D(N1073), .CK(clk), .Q(n3296) );
  DFFQX1 fft_d11_reg_26_ ( .D(N1105), .CK(clk), .Q(n3552) );
  DFFQX1 fft_d15_reg_26_ ( .D(stg_reg[26]), .CK(clk), .Q(n3680) );
  DFFQX1 fft_d3_reg_27_ ( .D(N1074), .CK(clk), .Q(n3295) );
  DFFQX1 fft_d7_reg_27_ ( .D(N1138), .CK(clk), .Q(n3423) );
  DFFQX1 fft_d11_reg_27_ ( .D(N1106), .CK(clk), .Q(n3551) );
  DFFQX1 fft_d15_reg_27_ ( .D(stg_reg[27]), .CK(clk), .Q(n3679) );
  DFFQX1 fft_d3_reg_28_ ( .D(N1075), .CK(clk), .Q(n3294) );
  DFFQX1 fft_d11_reg_28_ ( .D(N1107), .CK(clk), .Q(n3550) );
  DFFQX1 fft_d15_reg_28_ ( .D(stg_reg[28]), .CK(clk), .Q(n3678) );
  DFFQX1 fft_d3_reg_29_ ( .D(N1076), .CK(clk), .Q(n3293) );
  DFFQX1 fft_d7_reg_29_ ( .D(N1140), .CK(clk), .Q(n3421) );
  DFFQX1 fft_d15_reg_31_ ( .D(stg_reg[31]), .CK(clk), .Q(n3675) );
  DFFQX1 fft_d1_reg_6_ ( .D(N925), .CK(clk), .Q(n3252) );
  DFFQX1 fft_d1_reg_22_ ( .D(N941), .CK(clk), .Q(n3236) );
  DFFQX1 fft_d1_reg_5_ ( .D(N924), .CK(clk), .Q(n3253) );
  DFFQX1 fft_d1_reg_21_ ( .D(N940), .CK(clk), .Q(n3237) );
  DFFQX1 fft_d1_reg_4_ ( .D(N923), .CK(clk), .Q(n3254) );
  DFFQX1 fft_d1_reg_20_ ( .D(N939), .CK(clk), .Q(n3238) );
  DFFQX1 fft_d1_reg_3_ ( .D(N922), .CK(clk), .Q(n3255) );
  DFFQX1 fft_d1_reg_1_ ( .D(N920), .CK(clk), .Q(n3257) );
  DFFQX1 fft_d1_reg_17_ ( .D(N936), .CK(clk), .Q(n3241) );
  DFFQX1 fft_d1_reg_19_ ( .D(N938), .CK(clk), .Q(n3239) );
  DFFQX1 fft_d4_reg_0_ ( .D(N727), .CK(clk), .Q(n3354) );
  DFFQX1 fft_d12_reg_0_ ( .D(N759), .CK(clk), .Q(n3610) );
  DFFQX1 fft_d5_reg_1_ ( .D(N984), .CK(clk), .Q(n3385) );
  DFFQX1 fft_d9_reg_1_ ( .D(N952), .CK(clk), .Q(n3513) );
  DFFQX1 fft_d13_reg_1_ ( .D(N1016), .CK(clk), .Q(n3641) );
  DFFQX1 fft_d1_reg_2_ ( .D(N921), .CK(clk), .Q(n3256) );
  DFFQX1 fft_d5_reg_2_ ( .D(N985), .CK(clk), .Q(n3384) );
  DFFQX1 fft_d12_reg_2_ ( .D(N761), .CK(clk), .Q(n3608) );
  DFFQX1 fft_d5_reg_3_ ( .D(N986), .CK(clk), .Q(n3383) );
  DFFQX1 fft_d9_reg_3_ ( .D(N954), .CK(clk), .Q(n3511) );
  DFFQX1 fft_d13_reg_3_ ( .D(N1018), .CK(clk), .Q(n3639) );
  DFFQX1 fft_d5_reg_4_ ( .D(N987), .CK(clk), .Q(n3382) );
  DFFQX1 fft_d12_reg_4_ ( .D(N763), .CK(clk), .Q(n3606) );
  DFFQX1 fft_d5_reg_5_ ( .D(N988), .CK(clk), .Q(n3381) );
  DFFQX1 fft_d9_reg_5_ ( .D(N956), .CK(clk), .Q(n3509) );
  DFFQX1 fft_d13_reg_5_ ( .D(N1020), .CK(clk), .Q(n3637) );
  DFFQX1 fft_d5_reg_6_ ( .D(N989), .CK(clk), .Q(n3380) );
  DFFQX1 fft_d12_reg_6_ ( .D(N765), .CK(clk), .Q(n3604) );
  DFFQX1 fft_d1_reg_7_ ( .D(N926), .CK(clk), .Q(n3251) );
  DFFQX1 fft_d5_reg_7_ ( .D(N990), .CK(clk), .Q(n3379) );
  DFFQX1 fft_d9_reg_7_ ( .D(N958), .CK(clk), .Q(n3507) );
  DFFQX1 fft_d13_reg_7_ ( .D(N1022), .CK(clk), .Q(n3635) );
  DFFQX1 fft_d1_reg_8_ ( .D(N927), .CK(clk), .Q(n3250) );
  DFFQX1 fft_d5_reg_8_ ( .D(N991), .CK(clk), .Q(n3378) );
  DFFQX1 fft_d12_reg_8_ ( .D(N767), .CK(clk), .Q(n3602) );
  DFFQX1 fft_d1_reg_9_ ( .D(N928), .CK(clk), .Q(n3249) );
  DFFQX1 fft_d5_reg_9_ ( .D(N992), .CK(clk), .Q(n3377) );
  DFFQX1 fft_d9_reg_9_ ( .D(N960), .CK(clk), .Q(n3505) );
  DFFQX1 fft_d13_reg_9_ ( .D(N1024), .CK(clk), .Q(n3633) );
  DFFQX1 fft_d1_reg_10_ ( .D(N929), .CK(clk), .Q(n3248) );
  DFFQX1 fft_d5_reg_10_ ( .D(N993), .CK(clk), .Q(n3376) );
  DFFQX1 fft_d12_reg_10_ ( .D(N769), .CK(clk), .Q(n3600) );
  DFFQX1 fft_d1_reg_11_ ( .D(N930), .CK(clk), .Q(n3247) );
  DFFQX1 fft_d5_reg_11_ ( .D(N994), .CK(clk), .Q(n3375) );
  DFFQX1 fft_d9_reg_11_ ( .D(N962), .CK(clk), .Q(n3503) );
  DFFQX1 fft_d13_reg_11_ ( .D(N1026), .CK(clk), .Q(n3631) );
  DFFQX1 fft_d1_reg_12_ ( .D(N931), .CK(clk), .Q(n3246) );
  DFFQX1 fft_d5_reg_12_ ( .D(N995), .CK(clk), .Q(n3374) );
  DFFQX1 fft_d12_reg_12_ ( .D(N771), .CK(clk), .Q(n3598) );
  DFFQX1 fft_d1_reg_13_ ( .D(N932), .CK(clk), .Q(n3245) );
  DFFQX1 fft_d5_reg_13_ ( .D(N996), .CK(clk), .Q(n3373) );
  DFFQX1 fft_d9_reg_13_ ( .D(N964), .CK(clk), .Q(n3501) );
  DFFQX1 fft_d13_reg_13_ ( .D(N1028), .CK(clk), .Q(n3629) );
  DFFQX1 fft_d1_reg_14_ ( .D(N933), .CK(clk), .Q(n3244) );
  DFFQX1 fft_d5_reg_14_ ( .D(N997), .CK(clk), .Q(n3372) );
  DFFQX1 fft_d12_reg_14_ ( .D(N773), .CK(clk), .Q(n3596) );
  DFFQX1 fft_d5_reg_15_ ( .D(N998), .CK(clk), .Q(n3371) );
  DFFQX1 fft_d9_reg_15_ ( .D(N966), .CK(clk), .Q(n3499) );
  DFFQX1 fft_d13_reg_15_ ( .D(N1030), .CK(clk), .Q(n3627) );
  DFFQX1 fft_d1_reg_16_ ( .D(N935), .CK(clk), .Q(n3242) );
  DFFQX1 fft_d8_reg_16_ ( .D(N711), .CK(clk), .Q(n3466) );
  DFFQX1 fft_d13_reg_16_ ( .D(N1031), .CK(clk), .Q(n3626) );
  DFFQX1 fft_d5_reg_17_ ( .D(N1000), .CK(clk), .Q(n3369) );
  DFFQX1 fft_d9_reg_17_ ( .D(N968), .CK(clk), .Q(n3497) );
  DFFQX1 fft_d13_reg_17_ ( .D(N1032), .CK(clk), .Q(n3625) );
  DFFQX1 fft_d1_reg_18_ ( .D(N937), .CK(clk), .Q(n3240) );
  DFFQX1 fft_d8_reg_18_ ( .D(N713), .CK(clk), .Q(n3464) );
  DFFQX1 fft_d13_reg_18_ ( .D(N1033), .CK(clk), .Q(n3624) );
  DFFQX1 fft_d5_reg_19_ ( .D(N1002), .CK(clk), .Q(n3367) );
  DFFQX1 fft_d9_reg_19_ ( .D(N970), .CK(clk), .Q(n3495) );
  DFFQX1 fft_d13_reg_19_ ( .D(N1034), .CK(clk), .Q(n3623) );
  DFFQX1 fft_d8_reg_20_ ( .D(N715), .CK(clk), .Q(n3462) );
  DFFQX1 fft_d13_reg_20_ ( .D(N1035), .CK(clk), .Q(n3622) );
  DFFQX1 fft_d5_reg_21_ ( .D(N1004), .CK(clk), .Q(n3365) );
  DFFQX1 fft_d9_reg_21_ ( .D(N972), .CK(clk), .Q(n3493) );
  DFFQX1 fft_d13_reg_21_ ( .D(N1036), .CK(clk), .Q(n3621) );
  DFFQX1 fft_d8_reg_22_ ( .D(N717), .CK(clk), .Q(n3460) );
  DFFQX1 fft_d13_reg_22_ ( .D(N1037), .CK(clk), .Q(n3620) );
  DFFQX1 fft_d1_reg_23_ ( .D(N942), .CK(clk), .Q(n3235) );
  DFFQX1 fft_d5_reg_23_ ( .D(N1006), .CK(clk), .Q(n3363) );
  DFFQX1 fft_d9_reg_23_ ( .D(N974), .CK(clk), .Q(n3491) );
  DFFQX1 fft_d13_reg_23_ ( .D(N1038), .CK(clk), .Q(n3619) );
  DFFQX1 fft_d1_reg_24_ ( .D(N943), .CK(clk), .Q(n3234) );
  DFFQX1 fft_d8_reg_24_ ( .D(N719), .CK(clk), .Q(n3458) );
  DFFQX1 fft_d13_reg_24_ ( .D(N1039), .CK(clk), .Q(n3618) );
  DFFQX1 fft_d1_reg_25_ ( .D(N944), .CK(clk), .Q(n3233) );
  DFFQX1 fft_d5_reg_25_ ( .D(N1008), .CK(clk), .Q(n3361) );
  DFFQX1 fft_d9_reg_25_ ( .D(N976), .CK(clk), .Q(n3489) );
  DFFQX1 fft_d13_reg_25_ ( .D(N1040), .CK(clk), .Q(n3617) );
  DFFQX1 fft_d1_reg_26_ ( .D(N945), .CK(clk), .Q(n3232) );
  DFFQX1 fft_d8_reg_26_ ( .D(N721), .CK(clk), .Q(n3456) );
  DFFQX1 fft_d13_reg_26_ ( .D(N1041), .CK(clk), .Q(n3616) );
  DFFQX1 fft_d1_reg_27_ ( .D(N946), .CK(clk), .Q(n3231) );
  DFFQX1 fft_d5_reg_27_ ( .D(N1010), .CK(clk), .Q(n3359) );
  DFFQX1 fft_d9_reg_27_ ( .D(N978), .CK(clk), .Q(n3487) );
  DFFQX1 fft_d13_reg_27_ ( .D(N1042), .CK(clk), .Q(n3615) );
  DFFQX1 fft_d1_reg_28_ ( .D(N947), .CK(clk), .Q(n3230) );
  DFFQX1 fft_d8_reg_28_ ( .D(N723), .CK(clk), .Q(n3454) );
  DFFQX1 fft_d13_reg_28_ ( .D(N1043), .CK(clk), .Q(n3614) );
  DFFQX1 fft_d1_reg_29_ ( .D(N948), .CK(clk), .Q(n3229) );
  DFFQX1 fft_d5_reg_29_ ( .D(N1012), .CK(clk), .Q(n3357) );
  DFFQX1 fft_d12_reg_29_ ( .D(N788), .CK(clk), .Q(n3581) );
  DFFQX1 fft_d4_reg_30_ ( .D(N757), .CK(clk), .Q(n3324) );
  DFFQX1 fft_d8_reg_30_ ( .D(N725), .CK(clk), .Q(n3452) );
  DFFQX1 fft_d12_reg_30_ ( .D(N789), .CK(clk), .Q(n3580) );
  DFFQX1 fft_d4_reg_31_ ( .D(N758), .CK(clk), .Q(n3323) );
  DFFQX1 fft_d8_reg_31_ ( .D(N726), .CK(clk), .Q(n3451) );
  DFFQX1 fft_d12_reg_31_ ( .D(N790), .CK(clk), .Q(n3579) );
  DFFQX1 fft_d0_reg_13_ ( .D(N676), .CK(clk), .Q(n3721) );
  DFFQX1 fft_d0_reg_29_ ( .D(N692), .CK(clk), .Q(n3709) );
  DFFQX1 fft_d0_reg_9_ ( .D(N672), .CK(clk), .Q(n3725) );
  DFFQX1 fft_d0_reg_11_ ( .D(N674), .CK(clk), .Q(n3723) );
  DFFQX1 fft_d0_reg_27_ ( .D(N690), .CK(clk), .Q(n3711) );
  DFFQX1 fft_d0_reg_14_ ( .D(N677), .CK(clk), .Q(n3720) );
  DFFQX1 fft_d0_reg_30_ ( .D(N693), .CK(clk), .Q(n3708) );
  DFFQX1 fft_d3_reg_0_ ( .D(N1047), .CK(clk), .Q(n3322) );
  DFFQX1 fft_d11_reg_0_ ( .D(N1079), .CK(clk), .Q(n3578) );
  DFFQX1 fft_d11_reg_2_ ( .D(N1081), .CK(clk), .Q(n3576) );
  DFFQX1 fft_d11_reg_4_ ( .D(N1083), .CK(clk), .Q(n3574) );
  DFFQX1 fft_d11_reg_6_ ( .D(N1085), .CK(clk), .Q(n3572) );
  DFFQX1 fft_d11_reg_8_ ( .D(N1087), .CK(clk), .Q(n3570) );
  DFFQX1 fft_d11_reg_10_ ( .D(N1089), .CK(clk), .Q(n3568) );
  DFFQX1 fft_d11_reg_12_ ( .D(N1091), .CK(clk), .Q(n3566) );
  DFFQX1 fft_d11_reg_14_ ( .D(N1093), .CK(clk), .Q(n3564) );
  DFFQX1 fft_d7_reg_16_ ( .D(N1127), .CK(clk), .Q(n3434) );
  DFFQX1 fft_d7_reg_18_ ( .D(N1129), .CK(clk), .Q(n3432) );
  DFFQX1 fft_d7_reg_20_ ( .D(N1131), .CK(clk), .Q(n3430) );
  DFFQX1 fft_d7_reg_22_ ( .D(N1133), .CK(clk), .Q(n3428) );
  DFFQX1 fft_d7_reg_24_ ( .D(N1135), .CK(clk), .Q(n3426) );
  DFFQX1 fft_d7_reg_26_ ( .D(N1137), .CK(clk), .Q(n3424) );
  DFFQX1 fft_d7_reg_28_ ( .D(N1139), .CK(clk), .Q(n3422) );
  DFFQX1 fft_d11_reg_29_ ( .D(N1108), .CK(clk), .Q(n3549) );
  DFFQX1 fft_d15_reg_29_ ( .D(stg_reg[29]), .CK(clk), .Q(n3677) );
  DFFQX1 fft_d3_reg_30_ ( .D(N1077), .CK(clk), .Q(n3292) );
  DFFQX1 fft_d7_reg_30_ ( .D(N1141), .CK(clk), .Q(n3420) );
  DFFQX1 fft_d11_reg_30_ ( .D(N1109), .CK(clk), .Q(n3548) );
  DFFQX1 fft_d15_reg_30_ ( .D(stg_reg[30]), .CK(clk), .Q(n3676) );
  DFFQX1 fft_d3_reg_31_ ( .D(N1078), .CK(clk), .Q(n3291) );
  DFFQX1 fft_d7_reg_31_ ( .D(N1142), .CK(clk), .Q(n3419) );
  DFFQX1 fft_d11_reg_31_ ( .D(N1110), .CK(clk), .Q(n3547) );
  DFFQX1 fft_d1_reg_0_ ( .D(N919), .CK(clk), .Q(n3258) );
  DFFQX1 fft_d5_reg_0_ ( .D(N983), .CK(clk), .Q(n3386) );
  DFFQX1 fft_d8_reg_0_ ( .D(N695), .CK(clk), .Q(n3482) );
  DFFQX1 fft_d13_reg_0_ ( .D(N1015), .CK(clk), .Q(n3642) );
  DFFQX1 fft_d4_reg_1_ ( .D(N728), .CK(clk), .Q(n3353) );
  DFFQX1 fft_d8_reg_1_ ( .D(N696), .CK(clk), .Q(n3481) );
  DFFQX1 fft_d12_reg_1_ ( .D(N760), .CK(clk), .Q(n3609) );
  DFFQX1 fft_d4_reg_2_ ( .D(N729), .CK(clk), .Q(n3352) );
  DFFQX1 fft_d8_reg_2_ ( .D(N697), .CK(clk), .Q(n3480) );
  DFFQX1 fft_d13_reg_2_ ( .D(N1017), .CK(clk), .Q(n3640) );
  DFFQX1 fft_d4_reg_3_ ( .D(N730), .CK(clk), .Q(n3351) );
  DFFQX1 fft_d8_reg_3_ ( .D(N698), .CK(clk), .Q(n3479) );
  DFFQX1 fft_d12_reg_3_ ( .D(N762), .CK(clk), .Q(n3607) );
  DFFQX1 fft_d4_reg_4_ ( .D(N731), .CK(clk), .Q(n3350) );
  DFFQX1 fft_d8_reg_4_ ( .D(N699), .CK(clk), .Q(n3478) );
  DFFQX1 fft_d13_reg_4_ ( .D(N1019), .CK(clk), .Q(n3638) );
  DFFQX1 fft_d4_reg_5_ ( .D(N732), .CK(clk), .Q(n3349) );
  DFFQX1 fft_d8_reg_5_ ( .D(N700), .CK(clk), .Q(n3477) );
  DFFQX1 fft_d12_reg_5_ ( .D(N764), .CK(clk), .Q(n3605) );
  DFFQX1 fft_d4_reg_6_ ( .D(N733), .CK(clk), .Q(n3348) );
  DFFQX1 fft_d8_reg_6_ ( .D(N701), .CK(clk), .Q(n3476) );
  DFFQX1 fft_d13_reg_6_ ( .D(N1021), .CK(clk), .Q(n3636) );
  DFFQX1 fft_d4_reg_7_ ( .D(N734), .CK(clk), .Q(n3347) );
  DFFQX1 fft_d8_reg_7_ ( .D(N702), .CK(clk), .Q(n3475) );
  DFFQX1 fft_d12_reg_7_ ( .D(N766), .CK(clk), .Q(n3603) );
  DFFQX1 fft_d4_reg_8_ ( .D(N735), .CK(clk), .Q(n3346) );
  DFFQX1 fft_d8_reg_8_ ( .D(N703), .CK(clk), .Q(n3474) );
  DFFQX1 fft_d13_reg_8_ ( .D(N1023), .CK(clk), .Q(n3634) );
  DFFQX1 fft_d4_reg_9_ ( .D(N736), .CK(clk), .Q(n3345) );
  DFFQX1 fft_d8_reg_9_ ( .D(N704), .CK(clk), .Q(n3473) );
  DFFQX1 fft_d12_reg_9_ ( .D(N768), .CK(clk), .Q(n3601) );
  DFFQX1 fft_d4_reg_10_ ( .D(N737), .CK(clk), .Q(n3344) );
  DFFQX1 fft_d8_reg_10_ ( .D(N705), .CK(clk), .Q(n3472) );
  DFFQX1 fft_d13_reg_10_ ( .D(N1025), .CK(clk), .Q(n3632) );
  DFFQX1 fft_d4_reg_11_ ( .D(N738), .CK(clk), .Q(n3343) );
  DFFQX1 fft_d8_reg_11_ ( .D(N706), .CK(clk), .Q(n3471) );
  DFFQX1 fft_d12_reg_11_ ( .D(N770), .CK(clk), .Q(n3599) );
  DFFQX1 fft_d4_reg_12_ ( .D(N739), .CK(clk), .Q(n3342) );
  DFFQX1 fft_d8_reg_12_ ( .D(N707), .CK(clk), .Q(n3470) );
  DFFQX1 fft_d13_reg_12_ ( .D(N1027), .CK(clk), .Q(n3630) );
  DFFQX1 fft_d4_reg_13_ ( .D(N740), .CK(clk), .Q(n3341) );
  DFFQX1 fft_d8_reg_13_ ( .D(N708), .CK(clk), .Q(n3469) );
  DFFQX1 fft_d12_reg_13_ ( .D(N772), .CK(clk), .Q(n3597) );
  DFFQX1 fft_d4_reg_14_ ( .D(N741), .CK(clk), .Q(n3340) );
  DFFQX1 fft_d8_reg_14_ ( .D(N709), .CK(clk), .Q(n3468) );
  DFFQX1 fft_d13_reg_14_ ( .D(N1029), .CK(clk), .Q(n3628) );
  DFFQX1 fft_d1_reg_15_ ( .D(N934), .CK(clk), .Q(n3243) );
  DFFQX1 fft_d4_reg_15_ ( .D(N742), .CK(clk), .Q(n3339) );
  DFFQX1 fft_d8_reg_15_ ( .D(N710), .CK(clk), .Q(n3467) );
  DFFQX1 fft_d12_reg_15_ ( .D(N774), .CK(clk), .Q(n3595) );
  DFFQX1 fft_d4_reg_16_ ( .D(N743), .CK(clk), .Q(n3338) );
  DFFQX1 fft_d9_reg_16_ ( .D(N967), .CK(clk), .Q(n3498) );
  DFFQX1 fft_d12_reg_16_ ( .D(N775), .CK(clk), .Q(n3594) );
  DFFQX1 fft_d4_reg_17_ ( .D(N744), .CK(clk), .Q(n3337) );
  DFFQX1 fft_d8_reg_17_ ( .D(N712), .CK(clk), .Q(n3465) );
  DFFQX1 fft_d12_reg_17_ ( .D(N776), .CK(clk), .Q(n3593) );
  DFFQX1 fft_d4_reg_18_ ( .D(N745), .CK(clk), .Q(n3336) );
  DFFQX1 fft_d9_reg_18_ ( .D(N969), .CK(clk), .Q(n3496) );
  DFFQX1 fft_d12_reg_18_ ( .D(N777), .CK(clk), .Q(n3592) );
  DFFQX1 fft_d4_reg_19_ ( .D(N746), .CK(clk), .Q(n3335) );
  DFFQX1 fft_d8_reg_19_ ( .D(N714), .CK(clk), .Q(n3463) );
  DFFQX1 fft_d12_reg_19_ ( .D(N778), .CK(clk), .Q(n3591) );
  DFFQX1 fft_d4_reg_20_ ( .D(N747), .CK(clk), .Q(n3334) );
  DFFQX1 fft_d9_reg_20_ ( .D(N971), .CK(clk), .Q(n3494) );
  DFFQX1 fft_d12_reg_20_ ( .D(N779), .CK(clk), .Q(n3590) );
  DFFQX1 fft_d4_reg_21_ ( .D(N748), .CK(clk), .Q(n3333) );
  DFFQX1 fft_d8_reg_21_ ( .D(N716), .CK(clk), .Q(n3461) );
  DFFQX1 fft_d12_reg_21_ ( .D(N780), .CK(clk), .Q(n3589) );
  DFFQX1 fft_d4_reg_22_ ( .D(N749), .CK(clk), .Q(n3332) );
  DFFQX1 fft_d9_reg_22_ ( .D(N973), .CK(clk), .Q(n3492) );
  DFFQX1 fft_d12_reg_22_ ( .D(N781), .CK(clk), .Q(n3588) );
  DFFQX1 fft_d4_reg_23_ ( .D(N750), .CK(clk), .Q(n3331) );
  DFFQX1 fft_d8_reg_23_ ( .D(N718), .CK(clk), .Q(n3459) );
  DFFQX1 fft_d12_reg_23_ ( .D(N782), .CK(clk), .Q(n3587) );
  DFFQX1 fft_d4_reg_24_ ( .D(N751), .CK(clk), .Q(n3330) );
  DFFQX1 fft_d9_reg_24_ ( .D(N975), .CK(clk), .Q(n3490) );
  DFFQX1 fft_d12_reg_24_ ( .D(N783), .CK(clk), .Q(n3586) );
  DFFQX1 fft_d4_reg_25_ ( .D(N752), .CK(clk), .Q(n3329) );
  DFFQX1 fft_d8_reg_25_ ( .D(N720), .CK(clk), .Q(n3457) );
  DFFQX1 fft_d12_reg_25_ ( .D(N784), .CK(clk), .Q(n3585) );
  DFFQX1 fft_d4_reg_26_ ( .D(N753), .CK(clk), .Q(n3328) );
  DFFQX1 fft_d9_reg_26_ ( .D(N977), .CK(clk), .Q(n3488) );
  DFFQX1 fft_d12_reg_26_ ( .D(N785), .CK(clk), .Q(n3584) );
  DFFQX1 fft_d4_reg_27_ ( .D(N754), .CK(clk), .Q(n3327) );
  DFFQX1 fft_d8_reg_27_ ( .D(N722), .CK(clk), .Q(n3455) );
  DFFQX1 fft_d12_reg_27_ ( .D(N786), .CK(clk), .Q(n3583) );
  DFFQX1 fft_d4_reg_28_ ( .D(N755), .CK(clk), .Q(n3326) );
  DFFQX1 fft_d9_reg_28_ ( .D(N979), .CK(clk), .Q(n3486) );
  DFFQX1 fft_d12_reg_28_ ( .D(N787), .CK(clk), .Q(n3582) );
  DFFQX1 fft_d4_reg_29_ ( .D(N756), .CK(clk), .Q(n3325) );
  DFFQX1 fft_d8_reg_29_ ( .D(N724), .CK(clk), .Q(n3453) );
  DFFQX1 fft_d13_reg_29_ ( .D(N1044), .CK(clk), .Q(n3613) );
  DFFQX1 fft_d5_reg_30_ ( .D(N1013), .CK(clk), .Q(n3356) );
  DFFQX1 fft_d9_reg_30_ ( .D(N981), .CK(clk), .Q(n3484) );
  DFFQX1 fft_d13_reg_30_ ( .D(N1045), .CK(clk), .Q(n3612) );
  DFFQX1 fft_d1_reg_31_ ( .D(N950), .CK(clk), .Q(n3227) );
  DFFQX1 fft_d5_reg_31_ ( .D(N1014), .CK(clk), .Q(n3355) );
  DFFQX1 fft_d9_reg_31_ ( .D(N982), .CK(clk), .Q(n3483) );
  DFFQX1 fft_d13_reg_31_ ( .D(N1046), .CK(clk), .Q(n3611) );
  DFFHQX4 fft_d0_reg_16_ ( .D(N679), .CK(clk), .Q(n3718) );
  MDFFHQX1 fft_d2_reg_1_ ( .D0(stg_reg[129]), .D1(fft_d3[1]), .S0(n10330), 
        .CK(clk), .Q(n3289) );
  MDFFHQX1 fft_d2_reg_3_ ( .D0(stg_reg[131]), .D1(fft_d3[3]), .S0(n10320), 
        .CK(clk), .Q(n3287) );
  MDFFHQX1 fft_d2_reg_5_ ( .D0(stg_reg[133]), .D1(fft_d3[5]), .S0(n10310), 
        .CK(clk), .Q(n3285) );
  MDFFHQX1 fft_d2_reg_7_ ( .D0(stg_reg[135]), .D1(fft_d3[7]), .S0(n10300), 
        .CK(clk), .Q(n3283) );
  MDFFHQX1 fft_d2_reg_9_ ( .D0(stg_reg[137]), .D1(fft_d3[9]), .S0(n10290), 
        .CK(clk), .Q(n3281) );
  MDFFHQX1 fft_d2_reg_11_ ( .D0(stg_reg[139]), .D1(fft_d3[11]), .S0(n10280), 
        .CK(clk), .Q(n3279) );
  MDFFHQX1 fft_d2_reg_13_ ( .D0(stg_reg[141]), .D1(fft_d3[13]), .S0(n10270), 
        .CK(clk), .Q(n3277) );
  MDFFHQX1 fft_d6_reg_15_ ( .D0(stg_reg[79]), .D1(fft_d7[15]), .S0(n10260), 
        .CK(clk), .Q(n3403) );
  MDFFHQX1 fft_d14_reg_16_ ( .D0(stg_reg[48]), .D1(fft_d15[16]), .S0(n10250), 
        .CK(clk), .Q(n3658) );
  MDFFHQX1 fft_d14_reg_18_ ( .D0(stg_reg[50]), .D1(fft_d15[18]), .S0(n10240), 
        .CK(clk), .Q(n3656) );
  MDFFHQX1 fft_d14_reg_20_ ( .D0(stg_reg[52]), .D1(fft_d15[20]), .S0(n10230), 
        .CK(clk), .Q(n3654) );
  MDFFHQX1 fft_d14_reg_22_ ( .D0(stg_reg[54]), .D1(fft_d15[22]), .S0(n10220), 
        .CK(clk), .Q(n3652) );
  MDFFHQX1 fft_d14_reg_24_ ( .D0(stg_reg[56]), .D1(fft_d15[24]), .S0(n10210), 
        .CK(clk), .Q(n3650) );
  MDFFHQX1 fft_d14_reg_26_ ( .D0(stg_reg[58]), .D1(fft_d15[26]), .S0(n10200), 
        .CK(clk), .Q(n3648) );
  MDFFHQX1 fft_d14_reg_28_ ( .D0(stg_reg[60]), .D1(fft_d15[28]), .S0(n10190), 
        .CK(clk), .Q(n3646) );
  DFFQX1 fft_d0_reg_10_ ( .D(N673), .CK(clk), .Q(n3724) );
  DFFQX1 fft_d0_reg_26_ ( .D(N689), .CK(clk), .Q(n3712) );
  DFFQX1 fft_d0_reg_12_ ( .D(N675), .CK(clk), .Q(n3722) );
  DFFQX1 fft_d0_reg_28_ ( .D(N691), .CK(clk), .Q(n3710) );
  DFFQX1 fft_d9_reg_0_ ( .D(N951), .CK(clk), .Q(n3514) );
  DFFQX1 fft_d9_reg_2_ ( .D(N953), .CK(clk), .Q(n3512) );
  DFFQX1 fft_d9_reg_4_ ( .D(N955), .CK(clk), .Q(n3510) );
  DFFQX1 fft_d9_reg_6_ ( .D(N957), .CK(clk), .Q(n3508) );
  DFFQX1 fft_d9_reg_8_ ( .D(N959), .CK(clk), .Q(n3506) );
  DFFQX1 fft_d9_reg_10_ ( .D(N961), .CK(clk), .Q(n3504) );
  DFFQX1 fft_d9_reg_12_ ( .D(N963), .CK(clk), .Q(n3502) );
  DFFQX1 fft_d9_reg_14_ ( .D(N965), .CK(clk), .Q(n3500) );
  DFFQX1 fft_d5_reg_16_ ( .D(N999), .CK(clk), .Q(n3370) );
  DFFQX1 fft_d5_reg_18_ ( .D(N1001), .CK(clk), .Q(n3368) );
  DFFQX1 fft_d5_reg_20_ ( .D(N1003), .CK(clk), .Q(n3366) );
  DFFQX1 fft_d5_reg_22_ ( .D(N1005), .CK(clk), .Q(n3364) );
  DFFQX1 fft_d5_reg_24_ ( .D(N1007), .CK(clk), .Q(n3362) );
  DFFQX1 fft_d5_reg_26_ ( .D(N1009), .CK(clk), .Q(n3360) );
  DFFQX1 fft_d5_reg_28_ ( .D(N1011), .CK(clk), .Q(n3358) );
  DFFQX1 fft_d9_reg_29_ ( .D(N980), .CK(clk), .Q(n3485) );
  DFFQX1 fft_d1_reg_30_ ( .D(N949), .CK(clk), .Q(n3228) );
  DFFHQX4 fft_d0_reg_0_ ( .D(N663), .CK(clk), .Q(n3730) );
  MDFFHQX1 fft_d6_reg_0_ ( .D0(stg_reg[64]), .D1(fft_d7[0]), .S0(n10230), .CK(
        clk), .Q(n3418) );
  MDFFHQX1 fft_d14_reg_0_ ( .D0(stg_reg[32]), .D1(fft_d15[0]), .S0(n10330), 
        .CK(clk), .Q(n3674) );
  MDFFHQX1 fft_d14_reg_2_ ( .D0(stg_reg[34]), .D1(fft_d15[2]), .S0(n10320), 
        .CK(clk), .Q(n3672) );
  MDFFHQX1 fft_d14_reg_4_ ( .D0(stg_reg[36]), .D1(fft_d15[4]), .S0(n10310), 
        .CK(clk), .Q(n3670) );
  MDFFHQX1 fft_d14_reg_6_ ( .D0(stg_reg[38]), .D1(fft_d15[6]), .S0(n10300), 
        .CK(clk), .Q(n3668) );
  MDFFHQX1 fft_d14_reg_8_ ( .D0(stg_reg[40]), .D1(fft_d15[8]), .S0(n10290), 
        .CK(clk), .Q(n3666) );
  MDFFHQX1 fft_d14_reg_10_ ( .D0(stg_reg[42]), .D1(fft_d15[10]), .S0(n10280), 
        .CK(clk), .Q(n3664) );
  MDFFHQX1 fft_d14_reg_12_ ( .D0(stg_reg[44]), .D1(fft_d15[12]), .S0(n10270), 
        .CK(clk), .Q(n3662) );
  MDFFHQX1 fft_d14_reg_14_ ( .D0(stg_reg[46]), .D1(fft_d15[14]), .S0(n10260), 
        .CK(clk), .Q(n3660) );
  MDFFHQX1 fft_d10_reg_16_ ( .D0(stg_reg[112]), .D1(fft_d11[16]), .S0(n10250), 
        .CK(clk), .Q(n3530) );
  MDFFHQX1 fft_d10_reg_18_ ( .D0(stg_reg[114]), .D1(fft_d11[18]), .S0(n10240), 
        .CK(clk), .Q(n3528) );
  DFFQX1 stg_reg_reg_5__18_ ( .D(n2017), .CK(clk), .Q(stg_reg[114]) );
  MDFFHQX1 fft_d10_reg_20_ ( .D0(stg_reg[116]), .D1(fft_d11[20]), .S0(n10230), 
        .CK(clk), .Q(n3526) );
  MDFFHQX1 fft_d10_reg_22_ ( .D0(stg_reg[118]), .D1(fft_d11[22]), .S0(n10220), 
        .CK(clk), .Q(n3524) );
  MDFFHQX1 fft_d10_reg_24_ ( .D0(stg_reg[120]), .D1(fft_d11[24]), .S0(n10210), 
        .CK(clk), .Q(n3522) );
  MDFFHQX1 fft_d10_reg_26_ ( .D0(stg_reg[122]), .D1(fft_d11[26]), .S0(n10200), 
        .CK(clk), .Q(n3520) );
  MDFFHQX1 fft_d10_reg_28_ ( .D0(stg_reg[124]), .D1(fft_d11[28]), .S0(n10190), 
        .CK(clk), .Q(n3518) );
  MDFFHQX1 fft_d6_reg_1_ ( .D0(stg_reg[65]), .D1(fft_d7[1]), .S0(n10330), .CK(
        clk), .Q(n3417) );
  DFFQX1 stg_reg_reg_6__1_ ( .D(n1938), .CK(clk), .Q(stg_reg[65]) );
  MDFFHQX1 fft_d6_reg_3_ ( .D0(stg_reg[67]), .D1(fft_d7[3]), .S0(n10320), .CK(
        clk), .Q(n3415) );
  DFFQX1 stg_reg_reg_6__3_ ( .D(n1936), .CK(clk), .Q(stg_reg[67]) );
  MDFFHQX1 fft_d6_reg_5_ ( .D0(stg_reg[69]), .D1(fft_d7[5]), .S0(n10310), .CK(
        clk), .Q(n3413) );
  MDFFHQX1 fft_d6_reg_7_ ( .D0(stg_reg[71]), .D1(fft_d7[7]), .S0(n10300), .CK(
        clk), .Q(n3411) );
  MDFFHQX1 fft_d6_reg_9_ ( .D0(stg_reg[73]), .D1(fft_d7[9]), .S0(n10290), .CK(
        clk), .Q(n3409) );
  MDFFHQX1 fft_d6_reg_11_ ( .D0(stg_reg[75]), .D1(fft_d7[11]), .S0(n10280), 
        .CK(clk), .Q(n3407) );
  MDFFHQX1 fft_d6_reg_13_ ( .D0(stg_reg[77]), .D1(fft_d7[13]), .S0(n10270), 
        .CK(clk), .Q(n3405) );
  MDFFHQX1 fft_d2_reg_15_ ( .D0(stg_reg[143]), .D1(fft_d3[15]), .S0(n10260), 
        .CK(clk), .Q(n3275) );
  MDFFHQX1 fft_d2_reg_17_ ( .D0(stg_reg[145]), .D1(fft_d3[17]), .S0(n10250), 
        .CK(clk), .Q(n3273) );
  MDFFHQX1 fft_d2_reg_19_ ( .D0(stg_reg[147]), .D1(fft_d3[19]), .S0(n10240), 
        .CK(clk), .Q(n3271) );
  MDFFHQX1 fft_d2_reg_21_ ( .D0(stg_reg[149]), .D1(fft_d3[21]), .S0(n10230), 
        .CK(clk), .Q(n3269) );
  MDFFHQX1 fft_d2_reg_23_ ( .D0(stg_reg[151]), .D1(fft_d3[23]), .S0(n10220), 
        .CK(clk), .Q(n3267) );
  MDFFHQX1 fft_d2_reg_25_ ( .D0(stg_reg[153]), .D1(fft_d3[25]), .S0(n10210), 
        .CK(clk), .Q(n3265) );
  MDFFHQX1 fft_d2_reg_27_ ( .D0(stg_reg[155]), .D1(fft_d3[27]), .S0(n10200), 
        .CK(clk), .Q(n3263) );
  MDFFHQX1 fft_d2_reg_29_ ( .D0(stg_reg[157]), .D1(fft_d3[29]), .S0(n10190), 
        .CK(clk), .Q(n3261) );
  MDFFHQX1 fft_d10_reg_1_ ( .D0(stg_reg[97]), .D1(fft_d11[1]), .S0(n10330), 
        .CK(clk), .Q(n3545) );
  DFFQX1 stg_reg_reg_5__1_ ( .D(n2034), .CK(clk), .Q(stg_reg[97]) );
  MDFFHQX1 fft_d10_reg_3_ ( .D0(stg_reg[99]), .D1(fft_d11[3]), .S0(n10320), 
        .CK(clk), .Q(n3543) );
  DFFQX1 stg_reg_reg_5__3_ ( .D(n2032), .CK(clk), .Q(stg_reg[99]) );
  MDFFHQX1 fft_d10_reg_5_ ( .D0(stg_reg[101]), .D1(fft_d11[5]), .S0(n10310), 
        .CK(clk), .Q(n3541) );
  MDFFHQX1 fft_d10_reg_7_ ( .D0(stg_reg[103]), .D1(fft_d11[7]), .S0(n10300), 
        .CK(clk), .Q(n3539) );
  MDFFHQX1 fft_d10_reg_9_ ( .D0(stg_reg[105]), .D1(fft_d11[9]), .S0(n10290), 
        .CK(clk), .Q(n3537) );
  MDFFHQX1 fft_d10_reg_11_ ( .D0(stg_reg[107]), .D1(fft_d11[11]), .S0(n10280), 
        .CK(clk), .Q(n3535) );
  MDFFHQX1 fft_d10_reg_13_ ( .D0(stg_reg[109]), .D1(fft_d11[13]), .S0(n10270), 
        .CK(clk), .Q(n3533) );
  MDFFHQX1 fft_d10_reg_15_ ( .D0(stg_reg[111]), .D1(fft_d11[15]), .S0(n10260), 
        .CK(clk), .Q(n3531) );
  MDFFHQX1 fft_d6_reg_17_ ( .D0(stg_reg[81]), .D1(fft_d7[17]), .S0(n10250), 
        .CK(clk), .Q(n3401) );
  DFFQX1 stg_reg_reg_6__17_ ( .D(n1922), .CK(clk), .Q(stg_reg[81]) );
  MDFFHQX1 fft_d6_reg_19_ ( .D0(stg_reg[83]), .D1(fft_d7[19]), .S0(n10240), 
        .CK(clk), .Q(n3399) );
  DFFQX1 stg_reg_reg_6__19_ ( .D(n1920), .CK(clk), .Q(stg_reg[83]) );
  MDFFHQX1 fft_d6_reg_21_ ( .D0(stg_reg[85]), .D1(fft_d7[21]), .S0(n10230), 
        .CK(clk), .Q(n3397) );
  MDFFHQX1 fft_d6_reg_23_ ( .D0(stg_reg[87]), .D1(fft_d7[23]), .S0(n10220), 
        .CK(clk), .Q(n3395) );
  MDFFHQX1 fft_d6_reg_25_ ( .D0(stg_reg[89]), .D1(fft_d7[25]), .S0(n10210), 
        .CK(clk), .Q(n3393) );
  DFFQXL stg_reg_reg_6__25_ ( .D(n1914), .CK(clk), .Q(stg_reg[89]) );
  MDFFHQX1 fft_d6_reg_27_ ( .D0(stg_reg[91]), .D1(fft_d7[27]), .S0(n10200), 
        .CK(clk), .Q(n3391) );
  MDFFHQX1 fft_d6_reg_29_ ( .D0(stg_reg[93]), .D1(fft_d7[29]), .S0(n10190), 
        .CK(clk), .Q(n3389) );
  MDFFHQX1 fft_d14_reg_1_ ( .D0(stg_reg[33]), .D1(fft_d15[1]), .S0(n10330), 
        .CK(clk), .Q(n3673) );
  DFFQX1 stg_reg_reg_7__1_ ( .D(n1843), .CK(clk), .Q(stg_reg[33]) );
  MDFFHQX1 fft_d14_reg_3_ ( .D0(stg_reg[35]), .D1(fft_d15[3]), .S0(n10320), 
        .CK(clk), .Q(n3671) );
  DFFQX1 stg_reg_reg_7__3_ ( .D(n1841), .CK(clk), .Q(stg_reg[35]) );
  MDFFHQX1 fft_d14_reg_5_ ( .D0(stg_reg[37]), .D1(fft_d15[5]), .S0(n10310), 
        .CK(clk), .Q(n3669) );
  MDFFHQX1 fft_d14_reg_7_ ( .D0(stg_reg[39]), .D1(fft_d15[7]), .S0(n10300), 
        .CK(clk), .Q(n3667) );
  MDFFHQX1 fft_d14_reg_9_ ( .D0(stg_reg[41]), .D1(fft_d15[9]), .S0(n10290), 
        .CK(clk), .Q(n3665) );
  MDFFHQX1 fft_d14_reg_11_ ( .D0(stg_reg[43]), .D1(fft_d15[11]), .S0(n10280), 
        .CK(clk), .Q(n3663) );
  MDFFHQX1 fft_d14_reg_13_ ( .D0(stg_reg[45]), .D1(fft_d15[13]), .S0(n10270), 
        .CK(clk), .Q(n3661) );
  MDFFHQX1 fft_d14_reg_15_ ( .D0(stg_reg[47]), .D1(fft_d15[15]), .S0(n10260), 
        .CK(clk), .Q(n3659) );
  MDFFHQX1 fft_d10_reg_17_ ( .D0(stg_reg[113]), .D1(fft_d11[17]), .S0(n10250), 
        .CK(clk), .Q(n3529) );
  DFFQX1 stg_reg_reg_5__17_ ( .D(n2018), .CK(clk), .Q(stg_reg[113]) );
  MDFFHQX1 fft_d10_reg_19_ ( .D0(stg_reg[115]), .D1(fft_d11[19]), .S0(n10240), 
        .CK(clk), .Q(n3527) );
  DFFQX1 stg_reg_reg_5__19_ ( .D(n2016), .CK(clk), .Q(stg_reg[115]) );
  MDFFHQX1 fft_d10_reg_21_ ( .D0(stg_reg[117]), .D1(fft_d11[21]), .S0(n10230), 
        .CK(clk), .Q(n3525) );
  MDFFHQX1 fft_d10_reg_23_ ( .D0(stg_reg[119]), .D1(fft_d11[23]), .S0(n10220), 
        .CK(clk), .Q(n3523) );
  DFFQXL stg_reg_reg_5__23_ ( .D(n2012), .CK(clk), .Q(stg_reg[119]) );
  MDFFHQX1 fft_d10_reg_25_ ( .D0(stg_reg[121]), .D1(fft_d11[25]), .S0(n10210), 
        .CK(clk), .Q(n3521) );
  MDFFHQX1 fft_d10_reg_27_ ( .D0(stg_reg[123]), .D1(fft_d11[27]), .S0(n10200), 
        .CK(clk), .Q(n3519) );
  MDFFHQX1 fft_d2_reg_2_ ( .D0(stg_reg[130]), .D1(fft_d3[2]), .S0(n10330), 
        .CK(clk), .Q(n3288) );
  MDFFHQX1 fft_d2_reg_4_ ( .D0(stg_reg[132]), .D1(fft_d3[4]), .S0(n10320), 
        .CK(clk), .Q(n3286) );
  MDFFHQX1 fft_d2_reg_6_ ( .D0(stg_reg[134]), .D1(fft_d3[6]), .S0(n10310), 
        .CK(clk), .Q(n3284) );
  MDFFHQX1 fft_d2_reg_8_ ( .D0(stg_reg[136]), .D1(fft_d3[8]), .S0(n10300), 
        .CK(clk), .Q(n3282) );
  MDFFHQX1 fft_d2_reg_10_ ( .D0(stg_reg[138]), .D1(fft_d3[10]), .S0(n10290), 
        .CK(clk), .Q(n3280) );
  MDFFHQX1 fft_d2_reg_12_ ( .D0(stg_reg[140]), .D1(fft_d3[12]), .S0(n10280), 
        .CK(clk), .Q(n3278) );
  MDFFHQX1 fft_d2_reg_14_ ( .D0(stg_reg[142]), .D1(fft_d3[14]), .S0(n10270), 
        .CK(clk), .Q(n3276) );
  MDFFHQX1 fft_d2_reg_16_ ( .D0(stg_reg[144]), .D1(fft_d3[16]), .S0(n10260), 
        .CK(clk), .Q(n3274) );
  MDFFHQX1 fft_d14_reg_17_ ( .D0(stg_reg[49]), .D1(fft_d15[17]), .S0(n10250), 
        .CK(clk), .Q(n3657) );
  DFFQX1 stg_reg_reg_7__17_ ( .D(n1827), .CK(clk), .Q(stg_reg[49]) );
  MDFFHQX1 fft_d14_reg_19_ ( .D0(stg_reg[51]), .D1(fft_d15[19]), .S0(n10240), 
        .CK(clk), .Q(n3655) );
  DFFQX1 stg_reg_reg_7__19_ ( .D(n1825), .CK(clk), .Q(stg_reg[51]) );
  MDFFHQX1 fft_d14_reg_21_ ( .D0(stg_reg[53]), .D1(fft_d15[21]), .S0(n10230), 
        .CK(clk), .Q(n3653) );
  MDFFHQX1 fft_d14_reg_23_ ( .D0(stg_reg[55]), .D1(fft_d15[23]), .S0(n10220), 
        .CK(clk), .Q(n3651) );
  MDFFHQX1 fft_d14_reg_25_ ( .D0(stg_reg[57]), .D1(fft_d15[25]), .S0(n10210), 
        .CK(clk), .Q(n3649) );
  DFFQXL stg_reg_reg_7__25_ ( .D(n1819), .CK(clk), .Q(stg_reg[57]) );
  MDFFHQX1 fft_d14_reg_27_ ( .D0(stg_reg[59]), .D1(fft_d15[27]), .S0(n10200), 
        .CK(clk), .Q(n3647) );
  MDFFHQX1 fft_d6_reg_2_ ( .D0(stg_reg[66]), .D1(fft_d7[2]), .S0(n10330), .CK(
        clk), .Q(n3416) );
  MDFFHQX1 fft_d6_reg_4_ ( .D0(stg_reg[68]), .D1(fft_d7[4]), .S0(n10320), .CK(
        clk), .Q(n3414) );
  MDFFHQX1 fft_d6_reg_6_ ( .D0(stg_reg[70]), .D1(fft_d7[6]), .S0(n10310), .CK(
        clk), .Q(n3412) );
  MDFFHQX1 fft_d6_reg_8_ ( .D0(stg_reg[72]), .D1(fft_d7[8]), .S0(n10300), .CK(
        clk), .Q(n3410) );
  MDFFHQX1 fft_d6_reg_10_ ( .D0(stg_reg[74]), .D1(fft_d7[10]), .S0(n10290), 
        .CK(clk), .Q(n3408) );
  MDFFHQX1 fft_d6_reg_12_ ( .D0(stg_reg[76]), .D1(fft_d7[12]), .S0(n10280), 
        .CK(clk), .Q(n3406) );
  MDFFHQX1 fft_d6_reg_14_ ( .D0(stg_reg[78]), .D1(fft_d7[14]), .S0(n10270), 
        .CK(clk), .Q(n3404) );
  MDFFHQX1 fft_d2_reg_18_ ( .D0(stg_reg[146]), .D1(fft_d3[18]), .S0(n10250), 
        .CK(clk), .Q(n3272) );
  MDFFHQX1 fft_d2_reg_20_ ( .D0(stg_reg[148]), .D1(fft_d3[20]), .S0(n10240), 
        .CK(clk), .Q(n3270) );
  MDFFHQX1 fft_d2_reg_22_ ( .D0(stg_reg[150]), .D1(fft_d3[22]), .S0(n10230), 
        .CK(clk), .Q(n3268) );
  MDFFHQX1 fft_d2_reg_24_ ( .D0(stg_reg[152]), .D1(fft_d3[24]), .S0(n10220), 
        .CK(clk), .Q(n3266) );
  MDFFHQX1 fft_d2_reg_26_ ( .D0(stg_reg[154]), .D1(fft_d3[26]), .S0(n10210), 
        .CK(clk), .Q(n3264) );
  MDFFHQX1 fft_d2_reg_28_ ( .D0(stg_reg[156]), .D1(fft_d3[28]), .S0(n10200), 
        .CK(clk), .Q(n3262) );
  MDFFHQX1 fft_d14_reg_31_ ( .D0(stg_reg[63]), .D1(fft_d15[31]), .S0(n10260), 
        .CK(clk), .Q(n3643) );
  DFFXL stg_reg_reg_10__6_ ( .D(n1997), .CK(clk), .Q(n1570), .QN(n3119) );
  DFFXL stg_reg_reg_11__7_ ( .D(n1900), .CK(clk), .Q(n1608), .QN(n2967) );
  DFFXL stg_reg_reg_9__7_ ( .D(n2092), .CK(clk), .Q(n1525), .QN(n2968) );
  DFFXL stg_reg_reg_14__23_ ( .D(n1948), .CK(clk), .Q(n1750), .QN(n2782) );
  DFFXL stg_reg_reg_13__23_ ( .D(n2044), .CK(clk), .Q(n1702), .QN(n2784) );
  DFFXL stg_reg_reg_11__24_ ( .D(n1883), .CK(clk), .Q(n1786), .QN(n2771) );
  DFFXL stg_reg_reg_14__24_ ( .D(n1947), .CK(clk), .Q(n1753), .QN(n2772) );
  DFFXL stg_reg_reg_13__24_ ( .D(n2043), .CK(clk), .Q(n1705), .QN(n2774) );
  DFFXL stg_reg_reg_9__24_ ( .D(n2075), .CK(clk), .Q(n1704), .QN(n2773) );
  DFFXL stg_reg_reg_14__8_ ( .D(n1963), .CK(clk), .Q(n1577), .QN(n3111) );
  DFFXL stg_reg_reg_13__8_ ( .D(n2059), .CK(clk), .Q(n1529), .QN(n2956) );
  DFFXL stg_reg_reg_14__9_ ( .D(n1962), .CK(clk), .Q(n1580), .QN(n3106) );
  DFFXL stg_reg_reg_13__9_ ( .D(n2058), .CK(clk), .Q(n1532), .QN(n2943) );
  DFFXL stg_reg_reg_11__25_ ( .D(n1882), .CK(clk), .Q(n1788), .QN(n2761) );
  DFFXL stg_reg_reg_10__25_ ( .D(n1978), .CK(clk), .Q(n1755), .QN(n1344) );
  DFFXL stg_reg_reg_11__8_ ( .D(n1899), .CK(clk), .Q(n1610), .QN(n2954) );
  DFFXL stg_reg_reg_10__8_ ( .D(n1995), .CK(clk), .Q(n1576), .QN(n3110) );
  DFFXL stg_reg_reg_14__25_ ( .D(n1946), .CK(clk), .Q(n1756), .QN(n2762) );
  DFFXL stg_reg_reg_13__25_ ( .D(n2042), .CK(clk), .Q(n1708), .QN(n2764) );
  DFFXL stg_reg_reg_9__25_ ( .D(n2074), .CK(clk), .Q(n1707), .QN(n2763) );
  DFFXL stg_reg_reg_11__26_ ( .D(n1881), .CK(clk), .Q(n1760), .QN(n2751) );
  DFFXL stg_reg_reg_10__26_ ( .D(n1977), .CK(clk), .Q(n1713), .QN(n1335) );
  DFFXL stg_reg_reg_9__8_ ( .D(n2091), .CK(clk), .Q(n1528), .QN(n2955) );
  DFFXL stg_reg_reg_14__26_ ( .D(n1945), .CK(clk), .Q(n1714), .QN(n2752) );
  DFFXL stg_reg_reg_13__26_ ( .D(n2041), .CK(clk), .Q(n1666), .QN(n2754) );
  DFFXL stg_reg_reg_9__26_ ( .D(n2073), .CK(clk), .Q(n1665), .QN(n2753) );
  DFFXL stg_reg_reg_10__9_ ( .D(n1994), .CK(clk), .Q(n1579), .QN(n3105) );
  DFFXL stg_reg_reg_14__10_ ( .D(n1961), .CK(clk), .Q(n1538), .QN(n3102) );
  DFFXL stg_reg_reg_13__10_ ( .D(n2057), .CK(clk), .Q(n1490), .QN(n2930) );
  DFFXL stg_reg_reg_11__9_ ( .D(n1898), .CK(clk), .Q(n1612), .QN(n2941) );
  DFFXL stg_reg_reg_9__9_ ( .D(n2090), .CK(clk), .Q(n1531), .QN(n2942) );
  DFFXL stg_reg_reg_11__10_ ( .D(n1897), .CK(clk), .Q(n1584), .QN(n2928) );
  DFFXL stg_reg_reg_10__10_ ( .D(n1993), .CK(clk), .Q(n1537), .QN(n3101) );
  DFFXL stg_reg_reg_9__10_ ( .D(n2089), .CK(clk), .Q(n1489), .QN(n2929) );
  DFFXL stg_reg_reg_14__11_ ( .D(n1960), .CK(clk), .Q(n1541), .QN(n3098) );
  DFFXL stg_reg_reg_13__11_ ( .D(n2056), .CK(clk), .Q(n1493), .QN(n2917) );
  DFFXL stg_reg_reg_10__27_ ( .D(n1976), .CK(clk), .Q(n1716), .QN(n1326) );
  DFFXL stg_reg_reg_11__27_ ( .D(n1880), .CK(clk), .Q(n1762), .QN(n2741) );
  DFFXL stg_reg_reg_14__27_ ( .D(n1944), .CK(clk), .Q(n1717), .QN(n2742) );
  DFFXL stg_reg_reg_13__27_ ( .D(n2040), .CK(clk), .Q(n1669), .QN(n2744) );
  DFFXL stg_reg_reg_9__27_ ( .D(n2072), .CK(clk), .Q(n1668), .QN(n2743) );
  DFFXL stg_reg_reg_11__28_ ( .D(n1879), .CK(clk), .Q(n1764), .QN(n2731) );
  DFFXL stg_reg_reg_10__28_ ( .D(n1975), .CK(clk), .Q(n1719), .QN(n1317) );
  DFFXL stg_reg_reg_14__12_ ( .D(n1959), .CK(clk), .Q(n1544), .QN(n3094) );
  DFFXL stg_reg_reg_13__12_ ( .D(n2055), .CK(clk), .Q(n1496), .QN(n2904) );
  DFFXL stg_reg_reg_14__28_ ( .D(n1943), .CK(clk), .Q(n1720), .QN(n2732) );
  DFFXL stg_reg_reg_13__28_ ( .D(n2039), .CK(clk), .Q(n1672), .QN(n2734) );
  DFFXL stg_reg_reg_9__28_ ( .D(n2071), .CK(clk), .Q(n1671), .QN(n2733) );
  DFFXL stg_reg_reg_11__11_ ( .D(n1896), .CK(clk), .Q(n1586), .QN(n2915) );
  DFFXL stg_reg_reg_10__11_ ( .D(n1992), .CK(clk), .Q(n1540), .QN(n3097) );
  DFFXL stg_reg_reg_9__11_ ( .D(n2088), .CK(clk), .Q(n1492), .QN(n2916) );
  DFFXL stg_reg_reg_10__29_ ( .D(n1974), .CK(clk), .Q(n1722), .QN(n1308) );
  DFFXL stg_reg_reg_11__29_ ( .D(n1878), .CK(clk), .Q(n1766), .QN(n2721) );
  DFFXL stg_reg_reg_14__29_ ( .D(n1942), .CK(clk), .Q(n1723), .QN(n2722) );
  DFFXL stg_reg_reg_13__29_ ( .D(n2038), .CK(clk), .Q(n1675), .QN(n2724) );
  DFFXL stg_reg_reg_9__29_ ( .D(n2070), .CK(clk), .Q(n1674), .QN(n2723) );
  DFFXL stg_reg_reg_11__12_ ( .D(n1895), .CK(clk), .Q(n1588), .QN(n2902) );
  DFFXL stg_reg_reg_10__12_ ( .D(n1991), .CK(clk), .Q(n1543), .QN(n3093) );
  DFFXL stg_reg_reg_9__12_ ( .D(n2087), .CK(clk), .Q(n1495), .QN(n2903) );
  DFFXL stg_reg_reg_14__13_ ( .D(n1958), .CK(clk), .Q(n1547), .QN(n3090) );
  DFFXL stg_reg_reg_13__13_ ( .D(n2054), .CK(clk), .Q(n1499), .QN(n2891) );
  DFFXL stg_reg_reg_11__30_ ( .D(n1877), .CK(clk), .Q(n1768), .QN(n2712) );
  DFFXL stg_reg_reg_10__30_ ( .D(n1973), .CK(clk), .Q(n1725), .QN(n1297) );
  DFFXL stg_reg_reg_14__30_ ( .D(n1941), .CK(clk), .Q(n1726), .QN(n2713) );
  DFFXL stg_reg_reg_13__30_ ( .D(n2037), .CK(clk), .Q(n1678), .QN(n2714) );
  DFFRX2 cnt_reg_1_ ( .D(N36), .CK(clk), .RN(n3149), .Q(n109), .QN(n1811) );
  DFFQX1 fft_d0_reg_24_ ( .D(N687), .CK(clk), .Q(n3714) );
  DFFQX1 fft_d0_reg_23_ ( .D(N686), .CK(clk), .Q(n3715) );
  DFFQX1 fft_d0_reg_7_ ( .D(N670), .CK(clk), .Q(n3727) );
  DFFQX2 fft_d0_reg_18_ ( .D(N681), .CK(clk), .Q(fft_d0[18]) );
  DFFQX2 fft_d0_reg_2_ ( .D(N665), .CK(clk), .Q(fft_d0[2]) );
  DFFQX1 stg_reg_reg_15__0_ ( .D(n2308), .CK(clk), .Q(stg_reg[0]) );
  DFFQX1 stg_reg_reg_15__2_ ( .D(n1874), .CK(clk), .Q(stg_reg[2]) );
  DFFQX1 stg_reg_reg_15__18_ ( .D(n1858), .CK(clk), .Q(stg_reg[18]) );
  DFFQX1 stg_reg_reg_15__1_ ( .D(n1875), .CK(clk), .Q(stg_reg[1]) );
  DFFQX1 stg_reg_reg_15__3_ ( .D(n1873), .CK(clk), .Q(stg_reg[3]) );
  DFFQX2 fft_d0_reg_17_ ( .D(N680), .CK(clk), .Q(fft_d0[17]) );
  DFFQX1 stg_reg_reg_15__17_ ( .D(n1859), .CK(clk), .Q(stg_reg[17]) );
  DFFHQX4 fft_d0_reg_1_ ( .D(N664), .CK(clk), .Q(fft_d0[1]) );
  DFFQX4 fft_d0_reg_19_ ( .D(N682), .CK(clk), .Q(n3717) );
  DFFQX2 fft_d0_reg_3_ ( .D(N666), .CK(clk), .Q(n3729) );
  DFFHQX4 fft_d0_reg_20_ ( .D(N683), .CK(clk), .Q(fft_d0[20]) );
  DFFQX4 fft_d0_reg_4_ ( .D(N667), .CK(clk), .Q(fft_d0[4]) );
  DFFQX2 fft_d0_reg_22_ ( .D(N685), .CK(clk), .Q(n3716) );
  DFFQX2 fft_d0_reg_6_ ( .D(N669), .CK(clk), .Q(n3728) );
  DFFQX2 fft_d0_reg_21_ ( .D(N684), .CK(clk), .Q(fft_d0[21]) );
  DFFQX2 fft_d0_reg_5_ ( .D(N668), .CK(clk), .Q(fft_d0[5]) );
  DFFQX1 fft_d0_reg_8_ ( .D(N671), .CK(clk), .Q(n3726) );
  DFFQX1 fft_d0_reg_25_ ( .D(N688), .CK(clk), .Q(n3713) );
  DFFQX1 stg_reg_reg_15__29_ ( .D(n1847), .CK(clk), .Q(stg_reg[29]) );
  BUFX4 U3 ( .A(n9810), .Y(n9800) );
  CLKBUFX3 U4 ( .A(n3723), .Y(fft_d0[11]) );
  NAND4X2 U21 ( .A(n3014), .B(n3013), .C(n3012), .D(n3011), .Y(mul_1_in[4]) );
  OAI221X1 U22 ( .A0(n202), .A1(n1425), .B0(n77), .B1(n3071), .C0(n1423), .Y(
        n2004) );
  OAI221X4 U23 ( .A0(n9310), .A1(n3070), .B0(n9260), .B1(n3071), .C0(n1286), 
        .Y(n1940) );
  OAI221X4 U24 ( .A0(n51), .A1(n1425), .B0(n197), .B1(n3071), .C0(n1422), .Y(
        n2068) );
  OAI221X4 U49 ( .A0(n9310), .A1(n1425), .B0(n50), .B1(n3071), .C0(n1419), .Y(
        n2036) );
  INVX6 U50 ( .A(mul_o_sub[31]), .Y(n3071) );
  OAI221X2 U51 ( .A0(n9330), .A1(n2467), .B0(n854), .B1(n2869), .C0(n2464), 
        .Y(n1861) );
  OAI221X2 U52 ( .A0(n9330), .A1(n2566), .B0(n106), .B1(n2715), .C0(n2562), 
        .Y(n1846) );
  AOI2BB1X4 U53 ( .A0N(n2711), .A1N(n852), .B0(n822), .Y(n2562) );
  BUFX6 U54 ( .A(n3713), .Y(fft_d0[25]) );
  BUFX16 U55 ( .A(n7240), .Y(n17) );
  CLKBUFX2 U56 ( .A(n7240), .Y(n18) );
  BUFX20 U57 ( .A(n17), .Y(n19) );
  BUFX6 U58 ( .A(n17), .Y(n20) );
  CLKBUFX8 U59 ( .A(n17), .Y(n45) );
  CLKBUFX6 U60 ( .A(n17), .Y(n46) );
  CLKBUFX6 U61 ( .A(n17), .Y(n47) );
  BUFX12 U62 ( .A(n18), .Y(n48) );
  BUFX12 U63 ( .A(n18), .Y(n49) );
  BUFX12 U64 ( .A(n18), .Y(n50) );
  BUFX12 U65 ( .A(n18), .Y(n51) );
  BUFX12 U66 ( .A(n18), .Y(n52) );
  NAND2X1 U67 ( .A(n10430), .B(n109), .Y(n7240) );
  CLKINVX1 U68 ( .A(n9560), .Y(n53) );
  CLKINVX1 U69 ( .A(n53), .Y(n54) );
  CLKINVX1 U70 ( .A(n9550), .Y(n55) );
  CLKINVX1 U71 ( .A(n55), .Y(n56) );
  CLKINVX1 U72 ( .A(n9520), .Y(n57) );
  CLKINVX1 U73 ( .A(n57), .Y(n58) );
  CLKINVX1 U74 ( .A(n9530), .Y(n59) );
  CLKINVX1 U75 ( .A(n59), .Y(n60) );
  CLKINVX1 U76 ( .A(n9510), .Y(n61) );
  CLKINVX1 U77 ( .A(n61), .Y(n62) );
  CLKINVX1 U78 ( .A(n9540), .Y(n63) );
  CLKINVX1 U79 ( .A(n63), .Y(n64) );
  CLKINVX1 U80 ( .A(n9500), .Y(n65) );
  CLKINVX1 U81 ( .A(n65), .Y(n66) );
  CLKINVX1 U82 ( .A(n9490), .Y(n67) );
  CLKINVX1 U83 ( .A(n67), .Y(n68) );
  CLKINVX1 U84 ( .A(n9480), .Y(n69) );
  CLKINVX1 U85 ( .A(n69), .Y(n70) );
  CLKINVX1 U86 ( .A(n175), .Y(n71) );
  CLKINVX1 U87 ( .A(n71), .Y(n72) );
  CLKINVX12 U88 ( .A(n3144), .Y(n73) );
  CLKINVX4 U89 ( .A(n3144), .Y(n74) );
  INVX20 U90 ( .A(n73), .Y(n75) );
  INVX8 U91 ( .A(n73), .Y(n76) );
  INVX6 U92 ( .A(n73), .Y(n77) );
  INVX4 U93 ( .A(n73), .Y(n78) );
  INVX4 U94 ( .A(n73), .Y(n79) );
  INVX8 U95 ( .A(n74), .Y(n80) );
  INVX8 U96 ( .A(n74), .Y(n81) );
  INVX8 U97 ( .A(n74), .Y(n82) );
  INVX8 U98 ( .A(n74), .Y(n83) );
  INVX8 U99 ( .A(n74), .Y(n84) );
  NAND2X2 U100 ( .A(n837), .B(n10350), .Y(n3144) );
  CLKINVX1 U101 ( .A(n9480), .Y(n211) );
  INVXL U102 ( .A(n3144), .Y(n9560) );
  INVXL U103 ( .A(n3144), .Y(n9550) );
  CLKBUFX3 U104 ( .A(n9560), .Y(n9520) );
  CLKBUFX3 U105 ( .A(n9550), .Y(n9530) );
  CLKBUFX3 U106 ( .A(n9550), .Y(n9540) );
  CLKINVX1 U107 ( .A(n211), .Y(n175) );
  BUFX6 U108 ( .A(n3725), .Y(fft_d0[9]) );
  OAI221X2 U109 ( .A0(n9340), .A1(n2558), .B0(n106), .B1(n3073), .C0(n2554), 
        .Y(n1845) );
  AOI2BB1X4 U110 ( .A0N(n3071), .A1N(n852), .B0(n104), .Y(n2554) );
  BUFX6 U111 ( .A(n3715), .Y(fft_d0[23]) );
  BUFX6 U112 ( .A(n3714), .Y(fft_d0[24]) );
  BUFX6 U113 ( .A(n3726), .Y(fft_d0[8]) );
  CLKBUFX20 U114 ( .A(n3718), .Y(fft_d0[16]) );
  CLKINVX4 U115 ( .A(n468), .Y(fft_d0[7]) );
  CLKINVX4 U116 ( .A(n341), .Y(fft_d0[3]) );
  CLKINVX6 U117 ( .A(n10420), .Y(n10430) );
  AOI222X1 U118 ( .A0(stg_reg[49]), .A1(n861), .B0(stg_reg[81]), .B1(n913), 
        .C0(n1731), .C1(n904), .Y(n2850) );
  OA22X2 U119 ( .A0(n76), .A1(n3023), .B0(n10460), .B1(n3022), .Y(n3024) );
  AOI222XL U120 ( .A0(stg_reg[41]), .A1(n861), .B0(n914), .B1(stg_reg[73]), 
        .C0(n905), .C1(n1579), .Y(n2949) );
  INVX3 U121 ( .A(n1810), .Y(n10370) );
  OAI221X1 U122 ( .A0(n9740), .A1(n1147), .B0(n47), .B1(n1146), .C0(n1145), 
        .Y(stg2_img_Wn[48]) );
  CLKINVX1 U123 ( .A(mul_2_Wn_8), .Y(n2865) );
  AOI222X1 U124 ( .A0(stg_reg[33]), .A1(n862), .B0(n914), .B1(stg_reg[65]), 
        .C0(n905), .C1(n1555), .Y(n3053) );
  AOI222XL U125 ( .A0(stg_reg[36]), .A1(n862), .B0(n914), .B1(stg_reg[68]), 
        .C0(n904), .C1(n1564), .Y(n3014) );
  CLKBUFX3 U126 ( .A(mul_0_Wn[14]), .Y(n88) );
  AOI222X1 U127 ( .A0(stg_reg[57]), .A1(n862), .B0(stg_reg[89]), .B1(n914), 
        .C0(n1755), .C1(n905), .Y(n2770) );
  AOI222XL U128 ( .A0(stg_reg[56]), .A1(n862), .B0(stg_reg[88]), .B1(n913), 
        .C0(n1752), .C1(n904), .Y(n2780) );
  AOI222X1 U129 ( .A0(stg_reg[32]), .A1(n861), .B0(n914), .B1(stg_reg[64]), 
        .C0(n905), .C1(n1534), .Y(n3067) );
  BUFX4 U130 ( .A(mul_2_in[1]), .Y(n212) );
  NAND4X2 U131 ( .A(n2830), .B(n2829), .C(n2828), .D(n2827), .Y(mul_2_in[3])
         );
  AOI222XL U132 ( .A0(stg_reg[51]), .A1(n862), .B0(stg_reg[83]), .B1(n913), 
        .C0(n1737), .C1(n904), .Y(n2830) );
  AOI222X1 U133 ( .A0(stg_reg[55]), .A1(n862), .B0(stg_reg[87]), .B1(n914), 
        .C0(n1749), .C1(n905), .Y(n2790) );
  CLKBUFX3 U134 ( .A(n2949), .Y(n178) );
  CLKBUFX3 U135 ( .A(n2962), .Y(n179) );
  NAND4X1 U136 ( .A(n2988), .B(n2987), .C(n2986), .D(n2985), .Y(mul_1_in[6])
         );
  AOI222XL U137 ( .A0(stg_reg[38]), .A1(n861), .B0(n914), .B1(stg_reg[70]), 
        .C0(n905), .C1(n1570), .Y(n2988) );
  NAND4X4 U138 ( .A(n2975), .B(n2974), .C(n2973), .D(n2972), .Y(mul_1_in[7])
         );
  AOI222X1 U139 ( .A0(stg_reg[39]), .A1(n861), .B0(n914), .B1(stg_reg[71]), 
        .C0(n905), .C1(n1573), .Y(n2975) );
  AOI222XL U140 ( .A0(stg_reg[52]), .A1(n862), .B0(stg_reg[84]), .B1(n913), 
        .C0(n1740), .C1(n904), .Y(n2820) );
  NAND2X4 U141 ( .A(n7300), .B(n10460), .Y(mul_0_Wn_19) );
  CLKBUFX3 U142 ( .A(mul_0_Wn_1), .Y(n85) );
  NAND2X1 U143 ( .A(n2864), .B(n9670), .Y(mul_0_Wn_1) );
  NAND2X1 U144 ( .A(n3072), .B(n19), .Y(n10560) );
  INVX3 U145 ( .A(n85), .Y(n2861) );
  INVX3 U146 ( .A(n9710), .Y(n9670) );
  AND2X2 U147 ( .A(n867), .B(n9280), .Y(n7300) );
  CLKAND2X8 U148 ( .A(n909), .B(n75), .Y(n7320) );
  INVX3 U149 ( .A(n10560), .Y(n2864) );
  OAI221XL U150 ( .A0(n9800), .A1(n2845), .B0(n49), .B1(n2841), .C0(n2686), 
        .Y(stg2_real_Wn[1]) );
  OAI221X1 U151 ( .A0(n9780), .A1(n3061), .B0(n52), .B1(n3060), .C0(n2463), 
        .Y(stg2_img_Wn[32]) );
  OAI221X1 U152 ( .A0(n9750), .A1(n1283), .B0(n52), .B1(n1282), .C0(n1281), 
        .Y(stg2_real_Wn[48]) );
  AND2X2 U153 ( .A(n1811), .B(n838), .Y(n837) );
  BUFX16 U154 ( .A(n9250), .Y(n9280) );
  CLKBUFX3 U155 ( .A(n3072), .Y(n9210) );
  INVX4 U156 ( .A(n840), .Y(n3072) );
  CLKINVX1 U157 ( .A(stg_reg[119]), .Y(n2786) );
  CLKINVX1 U158 ( .A(stg_reg[115]), .Y(n2826) );
  CLKINVX1 U159 ( .A(stg_reg[99]), .Y(n3023) );
  CLKINVX1 U160 ( .A(stg_reg[114]), .Y(n2836) );
  CLKINVX1 U161 ( .A(stg_reg[98]), .Y(n3036) );
  CLKINVX1 U162 ( .A(stg_reg[20]), .Y(n2815) );
  CLKINVX1 U163 ( .A(stg_reg[101]), .Y(n2997) );
  CLKINVX1 U164 ( .A(stg_reg[117]), .Y(n2806) );
  CLKINVX1 U165 ( .A(stg_reg[5]), .Y(n2996) );
  CLKINVX1 U166 ( .A(stg_reg[21]), .Y(n2805) );
  CLKINVX1 U167 ( .A(stg_reg[19]), .Y(n2825) );
  INVX3 U168 ( .A(mul_o_sub[30]), .Y(n2711) );
  INVX3 U169 ( .A(mul_o_add[30]), .Y(n2878) );
  CLKINVX1 U170 ( .A(stg_reg[17]), .Y(n2845) );
  CLKINVX1 U171 ( .A(stg_reg[105]), .Y(n2945) );
  CLKINVX1 U172 ( .A(stg_reg[121]), .Y(n2766) );
  CLKINVX1 U173 ( .A(stg_reg[106]), .Y(n2932) );
  CLKINVX1 U174 ( .A(stg_reg[107]), .Y(n2919) );
  CLKINVX1 U175 ( .A(stg_reg[124]), .Y(n2736) );
  CLKINVX1 U176 ( .A(stg_reg[3]), .Y(n3022) );
  CLKINVX1 U177 ( .A(stg_reg[23]), .Y(n2785) );
  CLKINVX1 U178 ( .A(stg_reg[9]), .Y(n2944) );
  CLKINVX1 U179 ( .A(stg_reg[1]), .Y(n3048) );
  CLKINVX1 U180 ( .A(stg_reg[25]), .Y(n2765) );
  CLKINVX1 U181 ( .A(stg_reg[8]), .Y(n2957) );
  CLKINVX1 U182 ( .A(stg_reg[18]), .Y(n2835) );
  CLKINVX1 U183 ( .A(stg_reg[2]), .Y(n3035) );
  CLKINVX1 U184 ( .A(stg_reg[24]), .Y(n2775) );
  CLKINVX1 U185 ( .A(stg_reg[22]), .Y(n2795) );
  CLKINVX1 U186 ( .A(stg_reg[10]), .Y(n2931) );
  CLKINVX1 U187 ( .A(stg_reg[11]), .Y(n2918) );
  CLKINVX1 U188 ( .A(stg_reg[28]), .Y(n2735) );
  INVX6 U189 ( .A(n192), .Y(n193) );
  CLKINVX1 U190 ( .A(n9570), .Y(n192) );
  INVX4 U191 ( .A(n198), .Y(n199) );
  CLKINVX1 U192 ( .A(stg_reg[103]), .Y(n2971) );
  CLKINVX1 U193 ( .A(stg_reg[7]), .Y(n2970) );
  CLKINVX1 U194 ( .A(n9580), .Y(n190) );
  CLKINVX1 U195 ( .A(n9600), .Y(n194) );
  CLKBUFX3 U196 ( .A(n9540), .Y(n9490) );
  CLKINVX1 U197 ( .A(n9610), .Y(n196) );
  CLKINVX1 U198 ( .A(n9640), .Y(n188) );
  INVX3 U199 ( .A(n9650), .Y(n186) );
  CLKINVX1 U200 ( .A(n3729), .Y(n341) );
  CLKINVX1 U201 ( .A(n3727), .Y(n468) );
  CLKINVX16 U202 ( .A(n339), .Y(fft_d0[19]) );
  INVX3 U203 ( .A(n3717), .Y(n339) );
  BUFX12 U204 ( .A(n3675), .Y(fft_d15[31]) );
  BUFX12 U205 ( .A(n3294), .Y(fft_d3[28]) );
  BUFX12 U206 ( .A(n3296), .Y(fft_d3[26]) );
  BUFX12 U207 ( .A(n3298), .Y(fft_d3[24]) );
  BUFX12 U208 ( .A(n3300), .Y(fft_d3[22]) );
  BUFX12 U209 ( .A(n3302), .Y(fft_d3[20]) );
  BUFX12 U210 ( .A(n3304), .Y(fft_d3[18]) );
  BUFX12 U211 ( .A(n3436), .Y(fft_d7[14]) );
  BUFX12 U212 ( .A(n3438), .Y(fft_d7[12]) );
  BUFX12 U213 ( .A(n3440), .Y(fft_d7[10]) );
  BUFX12 U214 ( .A(n3442), .Y(fft_d7[8]) );
  BUFX12 U215 ( .A(n3444), .Y(fft_d7[6]) );
  BUFX12 U216 ( .A(n3446), .Y(fft_d7[4]) );
  BUFX12 U217 ( .A(n3448), .Y(fft_d7[2]) );
  BUFX12 U218 ( .A(n3679), .Y(fft_d15[27]) );
  BUFX12 U219 ( .A(n3681), .Y(fft_d15[25]) );
  BUFX12 U220 ( .A(n3683), .Y(fft_d15[23]) );
  BUFX12 U221 ( .A(n3685), .Y(fft_d15[21]) );
  BUFX12 U222 ( .A(n3687), .Y(fft_d15[19]) );
  BUFX12 U223 ( .A(n3689), .Y(fft_d15[17]) );
  BUFX12 U224 ( .A(n3306), .Y(fft_d3[16]) );
  BUFX12 U225 ( .A(n3308), .Y(fft_d3[14]) );
  BUFX12 U226 ( .A(n3310), .Y(fft_d3[12]) );
  BUFX12 U227 ( .A(n3312), .Y(fft_d3[10]) );
  BUFX12 U228 ( .A(n3314), .Y(fft_d3[8]) );
  BUFX12 U229 ( .A(n3316), .Y(fft_d3[6]) );
  BUFX12 U230 ( .A(n3318), .Y(fft_d3[4]) );
  BUFX12 U231 ( .A(n3320), .Y(fft_d3[2]) );
  BUFX12 U232 ( .A(n3551), .Y(fft_d11[27]) );
  BUFX12 U233 ( .A(n3553), .Y(fft_d11[25]) );
  BUFX12 U234 ( .A(n3555), .Y(fft_d11[23]) );
  BUFX12 U235 ( .A(n3557), .Y(fft_d11[21]) );
  BUFX12 U236 ( .A(n3559), .Y(fft_d11[19]) );
  BUFX12 U237 ( .A(n3561), .Y(fft_d11[17]) );
  BUFX12 U238 ( .A(n3691), .Y(fft_d15[15]) );
  BUFX12 U239 ( .A(n3693), .Y(fft_d15[13]) );
  BUFX12 U240 ( .A(n3695), .Y(fft_d15[11]) );
  BUFX12 U241 ( .A(n3697), .Y(fft_d15[9]) );
  BUFX12 U242 ( .A(n3699), .Y(fft_d15[7]) );
  BUFX12 U243 ( .A(n3701), .Y(fft_d15[5]) );
  BUFX12 U244 ( .A(n3703), .Y(fft_d15[3]) );
  BUFX12 U245 ( .A(n3705), .Y(fft_d15[1]) );
  BUFX12 U246 ( .A(n3421), .Y(fft_d7[29]) );
  BUFX12 U247 ( .A(n3423), .Y(fft_d7[27]) );
  BUFX12 U248 ( .A(n3425), .Y(fft_d7[25]) );
  BUFX12 U249 ( .A(n3427), .Y(fft_d7[23]) );
  BUFX12 U250 ( .A(n3429), .Y(fft_d7[21]) );
  BUFX12 U251 ( .A(n3431), .Y(fft_d7[19]) );
  BUFX12 U252 ( .A(n3433), .Y(fft_d7[17]) );
  BUFX12 U253 ( .A(n3563), .Y(fft_d11[15]) );
  BUFX12 U254 ( .A(n3565), .Y(fft_d11[13]) );
  BUFX12 U255 ( .A(n3567), .Y(fft_d11[11]) );
  BUFX12 U256 ( .A(n3569), .Y(fft_d11[9]) );
  BUFX12 U257 ( .A(n3571), .Y(fft_d11[7]) );
  BUFX12 U258 ( .A(n3573), .Y(fft_d11[5]) );
  BUFX12 U259 ( .A(n3575), .Y(fft_d11[3]) );
  BUFX12 U260 ( .A(n3577), .Y(fft_d11[1]) );
  BUFX12 U261 ( .A(n3293), .Y(fft_d3[29]) );
  BUFX12 U262 ( .A(n3295), .Y(fft_d3[27]) );
  BUFX12 U263 ( .A(n3297), .Y(fft_d3[25]) );
  BUFX12 U264 ( .A(n3299), .Y(fft_d3[23]) );
  BUFX12 U265 ( .A(n3301), .Y(fft_d3[21]) );
  BUFX12 U266 ( .A(n3303), .Y(fft_d3[19]) );
  BUFX12 U267 ( .A(n3305), .Y(fft_d3[17]) );
  BUFX12 U268 ( .A(n3307), .Y(fft_d3[15]) );
  BUFX12 U269 ( .A(n3437), .Y(fft_d7[13]) );
  BUFX12 U270 ( .A(n3439), .Y(fft_d7[11]) );
  BUFX12 U271 ( .A(n3441), .Y(fft_d7[9]) );
  BUFX12 U272 ( .A(n3443), .Y(fft_d7[7]) );
  BUFX12 U273 ( .A(n3445), .Y(fft_d7[5]) );
  BUFX12 U274 ( .A(n3447), .Y(fft_d7[3]) );
  BUFX12 U275 ( .A(n3449), .Y(fft_d7[1]) );
  BUFX12 U276 ( .A(n3550), .Y(fft_d11[28]) );
  BUFX12 U277 ( .A(n3552), .Y(fft_d11[26]) );
  BUFX12 U278 ( .A(n3554), .Y(fft_d11[24]) );
  BUFX12 U279 ( .A(n3556), .Y(fft_d11[22]) );
  BUFX12 U280 ( .A(n3558), .Y(fft_d11[20]) );
  BUFX12 U281 ( .A(n3560), .Y(fft_d11[18]) );
  BUFX12 U282 ( .A(n3562), .Y(fft_d11[16]) );
  BUFX12 U283 ( .A(n3692), .Y(fft_d15[14]) );
  BUFX12 U284 ( .A(n3694), .Y(fft_d15[12]) );
  BUFX12 U285 ( .A(n3696), .Y(fft_d15[10]) );
  BUFX12 U286 ( .A(n3698), .Y(fft_d15[8]) );
  BUFX12 U287 ( .A(n3700), .Y(fft_d15[6]) );
  BUFX12 U288 ( .A(n3702), .Y(fft_d15[4]) );
  BUFX12 U289 ( .A(n3704), .Y(fft_d15[2]) );
  BUFX12 U290 ( .A(n3706), .Y(fft_d15[0]) );
  BUFX12 U291 ( .A(n3450), .Y(fft_d7[0]) );
  BUFX12 U292 ( .A(n3678), .Y(fft_d15[28]) );
  BUFX12 U293 ( .A(n3680), .Y(fft_d15[26]) );
  BUFX12 U294 ( .A(n3682), .Y(fft_d15[24]) );
  BUFX12 U295 ( .A(n3684), .Y(fft_d15[22]) );
  BUFX12 U296 ( .A(n3686), .Y(fft_d15[20]) );
  BUFX12 U297 ( .A(n3688), .Y(fft_d15[18]) );
  BUFX12 U298 ( .A(n3690), .Y(fft_d15[16]) );
  BUFX12 U299 ( .A(n3435), .Y(fft_d7[15]) );
  BUFX12 U300 ( .A(n3309), .Y(fft_d3[13]) );
  BUFX12 U301 ( .A(n3311), .Y(fft_d3[11]) );
  BUFX12 U302 ( .A(n3313), .Y(fft_d3[9]) );
  BUFX12 U303 ( .A(n3315), .Y(fft_d3[7]) );
  BUFX12 U304 ( .A(n3317), .Y(fft_d3[5]) );
  BUFX12 U305 ( .A(n3319), .Y(fft_d3[3]) );
  BUFX12 U306 ( .A(n3321), .Y(fft_d3[1]) );
  OAI221X1 U307 ( .A0(n902), .A1(n150), .B0(n890), .B1(n2867), .C0(n2866), .Y(
        n1988) );
  OAI221X1 U308 ( .A0(n855), .A1(n111), .B0(n893), .B1(n2466), .C0(n2465), .Y(
        n1892) );
  NAND4X2 U309 ( .A(n2820), .B(n2819), .C(n2818), .D(n2817), .Y(mul_2_in[4])
         );
  NAND2X4 U310 ( .A(n2864), .B(n10440), .Y(mul_2_Wn_9) );
  CLKBUFX3 U311 ( .A(mul_0_Wn_2), .Y(n86) );
  BUFX4 U312 ( .A(mul_0_Wn_2), .Y(n87) );
  NAND2X1 U313 ( .A(n2864), .B(n2863), .Y(mul_0_Wn_2) );
  NAND2XL U314 ( .A(n7300), .B(n2861), .Y(mul_0_Wn[14]) );
  INVX3 U315 ( .A(n9720), .Y(n9690) );
  INVX8 U316 ( .A(n182), .Y(n183) );
  NAND2XL U317 ( .A(n850), .B(n185), .Y(n3142) );
  INVX4 U318 ( .A(n184), .Y(n185) );
  INVX6 U319 ( .A(n190), .Y(n191) );
  INVX2 U320 ( .A(n9710), .Y(n9680) );
  INVX4 U321 ( .A(n180), .Y(n181) );
  INVX3 U322 ( .A(n184), .Y(n200) );
  INVX6 U323 ( .A(n196), .Y(n197) );
  INVX4 U324 ( .A(n180), .Y(n203) );
  INVX3 U325 ( .A(n201), .Y(n202) );
  CLKINVX1 U326 ( .A(n9710), .Y(n9590) );
  INVX6 U327 ( .A(n188), .Y(n189) );
  INVX3 U328 ( .A(n9660), .Y(n198) );
  INVX6 U329 ( .A(n194), .Y(n195) );
  INVX8 U330 ( .A(n186), .Y(n187) );
  CLKINVX1 U331 ( .A(n9720), .Y(n9630) );
  INVX4 U332 ( .A(n206), .Y(n207) );
  INVX4 U333 ( .A(n915), .Y(n914) );
  CLKBUFX3 U334 ( .A(n7250), .Y(n863) );
  INVX3 U335 ( .A(n204), .Y(n205) );
  INVX8 U336 ( .A(n909), .Y(n904) );
  INVX6 U337 ( .A(n907), .Y(n905) );
  CLKBUFX6 U338 ( .A(n7260), .Y(n915) );
  NAND2X2 U339 ( .A(n791), .B(n10350), .Y(n7250) );
  INVX3 U340 ( .A(n9670), .Y(n201) );
  INVX3 U341 ( .A(n9690), .Y(n180) );
  BUFX6 U342 ( .A(n903), .Y(n909) );
  NAND2X2 U343 ( .A(n10530), .B(n10350), .Y(n7260) );
  NAND3BXL U344 ( .AN(n209), .B(n52), .C(n77), .Y(n3148) );
  INVX3 U345 ( .A(n9700), .Y(n184) );
  CLKBUFX3 U346 ( .A(n9540), .Y(n9480) );
  BUFX6 U347 ( .A(n3055), .Y(n903) );
  BUFX12 U348 ( .A(n9730), .Y(n9710) );
  INVX3 U349 ( .A(n9660), .Y(n204) );
  CLKBUFX2 U350 ( .A(n903), .Y(n906) );
  CLKBUFX3 U351 ( .A(n9730), .Y(n9720) );
  INVX3 U352 ( .A(n9680), .Y(n206) );
  AND2X2 U353 ( .A(stg2_real_14__15_), .B(n880), .Y(n103) );
  AND2X2 U354 ( .A(stg2_real_15__15_), .B(n884), .Y(n104) );
  AND2X2 U355 ( .A(n1300), .B(n10520), .Y(n106) );
  AND4XL U356 ( .A(n1287), .B(n187), .C(n9200), .D(n77), .Y(n107) );
  AND4XL U357 ( .A(n1301), .B(n7300), .C(n852), .D(n1300), .Y(n153) );
  BUFX2 U358 ( .A(n7250), .Y(n867) );
  AOI222XL U359 ( .A0(stg_reg[58]), .A1(n862), .B0(stg_reg[90]), .B1(n914), 
        .C0(n1713), .C1(n905), .Y(n2760) );
  AND2X2 U360 ( .A(stg2_real_13__15_), .B(n881), .Y(n120) );
  XNOR2X1 U361 ( .A(n3164), .B(n7850), .Y(n121) );
  XNOR2X1 U362 ( .A(n3163), .B(n7820), .Y(n122) );
  XNOR2X1 U363 ( .A(n3165), .B(n7880), .Y(n123) );
  XNOR2X1 U364 ( .A(n3162), .B(n7790), .Y(n129) );
  XNOR2X1 U365 ( .A(n3161), .B(n7760), .Y(n130) );
  XNOR2X1 U366 ( .A(n3160), .B(n7730), .Y(n131) );
  XNOR2X1 U367 ( .A(n3159), .B(n7700), .Y(n147) );
  XNOR2X1 U368 ( .A(n3158), .B(n7670), .Y(n148) );
  XNOR2X1 U369 ( .A(n3157), .B(n7520), .Y(n149) );
  CLKINVX1 U370 ( .A(n1285), .Y(n3079) );
  CLKINVX1 U371 ( .A(n1418), .Y(n2456) );
  CLKINVX1 U372 ( .A(n10590), .Y(n2460) );
  CLKINVX1 U373 ( .A(n10580), .Y(n2690) );
  CLKINVX1 U374 ( .A(n1421), .Y(n2458) );
  XNOR2X1 U375 ( .A(n3156), .B(n7640), .Y(n162) );
  XNOR2X1 U376 ( .A(n3155), .B(n7490), .Y(n163) );
  XNOR2X1 U377 ( .A(n3154), .B(n7610), .Y(n164) );
  AND2X2 U378 ( .A(stg2_real_14__0_), .B(n882), .Y(n165) );
  AND2X2 U379 ( .A(stg2_real_15__0_), .B(n886), .Y(n166) );
  AND2X2 U380 ( .A(stg2_real_13__0_), .B(n886), .Y(n167) );
  XNOR2X1 U381 ( .A(n3151), .B(n3150), .Y(n172) );
  XNOR2X1 U382 ( .A(n3153), .B(n7580), .Y(n173) );
  XNOR2X1 U383 ( .A(n3152), .B(n7550), .Y(n174) );
  NAND2X1 U384 ( .A(n10480), .B(n10350), .Y(n3082) );
  CLKINVX1 U385 ( .A(n1810), .Y(n10360) );
  INVX4 U386 ( .A(mul_2_Wn[13]), .Y(n10460) );
  NAND3BX1 U387 ( .AN(n176), .B(n1811), .C(n177), .Y(n10450) );
  CLKAND2X4 U388 ( .A(n10430), .B(n1811), .Y(n841) );
  AOI222X4 U389 ( .A0(stg_reg[34]), .A1(n862), .B0(n914), .B1(stg_reg[66]), 
        .C0(n904), .C1(n1558), .Y(n3040) );
  NAND2XL U390 ( .A(n837), .B(n10360), .Y(n2687) );
  BUFX2 U391 ( .A(n3072), .Y(n9220) );
  CLKBUFX3 U392 ( .A(n9220), .Y(n918) );
  CLKBUFX4 U393 ( .A(n9220), .Y(n917) );
  NAND4X2 U394 ( .A(n2760), .B(n2759), .C(n2758), .D(n2757), .Y(mul_2_in[10])
         );
  CLKINVX8 U395 ( .A(n9620), .Y(n182) );
  INVXL U396 ( .A(n839), .Y(n208) );
  INVX3 U397 ( .A(n208), .Y(n209) );
  BUFX4 U398 ( .A(n839), .Y(n9730) );
  INVX4 U399 ( .A(n198), .Y(n9620) );
  CLKINVX3 U400 ( .A(n201), .Y(n9700) );
  INVX2 U401 ( .A(n9720), .Y(n9650) );
  INVX1 U402 ( .A(n206), .Y(n9640) );
  INVXL U403 ( .A(n204), .Y(n9580) );
  INVXL U404 ( .A(n198), .Y(n9570) );
  INVXL U405 ( .A(n9710), .Y(n9600) );
  INVXL U406 ( .A(n9710), .Y(n9610) );
  INVX4 U407 ( .A(n9710), .Y(n9660) );
  NAND4X4 U408 ( .A(n3027), .B(n3026), .C(n3025), .D(n3024), .Y(mul_1_in[3])
         );
  AOI222X4 U409 ( .A0(stg_reg[35]), .A1(n861), .B0(n914), .B1(stg_reg[67]), 
        .C0(n905), .C1(n1561), .Y(n3027) );
  BUFX3 U410 ( .A(n3001), .Y(n210) );
  NAND2X4 U411 ( .A(n7320), .B(n2862), .Y(mul_2_Wn[14]) );
  INVX3 U412 ( .A(mul_0_Wn_19), .Y(n2862) );
  NAND4X4 U413 ( .A(n2730), .B(n2729), .C(n2728), .D(n2727), .Y(mul_2_in[13])
         );
  AOI222X4 U414 ( .A0(stg_reg[61]), .A1(n862), .B0(stg_reg[93]), .B1(n913), 
        .C0(n1722), .C1(n904), .Y(n2730) );
  NAND4X6 U415 ( .A(n2750), .B(n2749), .C(n2748), .D(n2747), .Y(mul_2_in[11])
         );
  AOI222X4 U416 ( .A0(stg_reg[59]), .A1(n862), .B0(stg_reg[91]), .B1(n914), 
        .C0(n1716), .C1(n905), .Y(n2750) );
  NAND4X4 U417 ( .A(n2810), .B(n2809), .C(n2808), .D(n2807), .Y(mul_2_in[5])
         );
  AOI222X4 U418 ( .A0(stg_reg[53]), .A1(n862), .B0(stg_reg[85]), .B1(n913), 
        .C0(n1743), .C1(n904), .Y(n2810) );
  AOI222X4 U419 ( .A0(stg_reg[50]), .A1(n861), .B0(stg_reg[82]), .B1(n913), 
        .C0(n1734), .C1(n904), .Y(n2840) );
  NAND3BX2 U420 ( .AN(n177), .B(n1810), .C(n176), .Y(n10420) );
  OA22X4 U421 ( .A0(n77), .A1(n3049), .B0(n10460), .B1(n3048), .Y(n3050) );
  INVX8 U422 ( .A(n10370), .Y(n10350) );
  NAND4X4 U423 ( .A(n3040), .B(n3039), .C(n3038), .D(n3037), .Y(mul_1_in[2])
         );
  NAND4X4 U424 ( .A(n2860), .B(n2859), .C(n2858), .D(n2857), .Y(mul_2_in[0])
         );
  AOI222X4 U425 ( .A0(stg_reg[48]), .A1(n861), .B0(stg_reg[80]), .B1(n913), 
        .C0(n1710), .C1(n904), .Y(n2860) );
  CLKBUFX2 U426 ( .A(n9560), .Y(n9510) );
  CLKBUFX2 U427 ( .A(n9520), .Y(n9500) );
  NAND4X4 U428 ( .A(n210), .B(n3000), .C(n2999), .D(n2998), .Y(mul_1_in[5]) );
  OAI221X2 U429 ( .A0(n848), .A1(n2868), .B0(n896), .B1(n2389), .C0(n2388), 
        .Y(n2084) );
  INVXL U430 ( .A(mul_2_Wn_9), .Y(n10470) );
  AND4X1 U431 ( .A(n1790), .B(n109), .C(n177), .D(n1810), .Y(n839) );
  INVX8 U432 ( .A(n916), .Y(n913) );
  NAND4X4 U433 ( .A(n2770), .B(n2769), .C(n2768), .D(n2767), .Y(mul_2_in[9])
         );
  NAND4X4 U434 ( .A(n2790), .B(n2789), .C(n2788), .D(n2787), .Y(mul_2_in[7])
         );
  NAND4X4 U435 ( .A(n2800), .B(n2799), .C(n2798), .D(n2797), .Y(mul_2_in[6])
         );
  OA22XL U436 ( .A0(n78), .A1(n2796), .B0(n10350), .B1(n2795), .Y(n2797) );
  AOI222X4 U437 ( .A0(stg_reg[54]), .A1(n862), .B0(stg_reg[86]), .B1(n913), 
        .C0(n1746), .C1(n904), .Y(n2800) );
  NAND4X4 U438 ( .A(n2840), .B(n2839), .C(n2838), .D(n2837), .Y(mul_2_in[2])
         );
  BUFX12 U439 ( .A(n3643), .Y(fft_d14[31]) );
  BUFX12 U440 ( .A(n3262), .Y(fft_d2[28]) );
  BUFX12 U441 ( .A(n3264), .Y(fft_d2[26]) );
  BUFX12 U442 ( .A(n3266), .Y(fft_d2[24]) );
  BUFX12 U443 ( .A(n3268), .Y(fft_d2[22]) );
  BUFX12 U444 ( .A(n3270), .Y(fft_d2[20]) );
  BUFX12 U445 ( .A(n3272), .Y(fft_d2[18]) );
  BUFX12 U446 ( .A(n3404), .Y(fft_d6[14]) );
  BUFX12 U447 ( .A(n3406), .Y(fft_d6[12]) );
  BUFX12 U448 ( .A(n3408), .Y(fft_d6[10]) );
  BUFX12 U449 ( .A(n3410), .Y(fft_d6[8]) );
  BUFX12 U450 ( .A(n3412), .Y(fft_d6[6]) );
  BUFX12 U451 ( .A(n3414), .Y(fft_d6[4]) );
  BUFX12 U452 ( .A(n3416), .Y(fft_d6[2]) );
  BUFX12 U453 ( .A(n3647), .Y(fft_d14[27]) );
  BUFX12 U454 ( .A(n3649), .Y(fft_d14[25]) );
  BUFX12 U455 ( .A(n3651), .Y(fft_d14[23]) );
  BUFX12 U456 ( .A(n3653), .Y(fft_d14[21]) );
  BUFX12 U457 ( .A(n3655), .Y(fft_d14[19]) );
  BUFX12 U458 ( .A(n3657), .Y(fft_d14[17]) );
  BUFX12 U459 ( .A(n3274), .Y(fft_d2[16]) );
  BUFX12 U460 ( .A(n3276), .Y(fft_d2[14]) );
  BUFX12 U461 ( .A(n3278), .Y(fft_d2[12]) );
  BUFX12 U462 ( .A(n3280), .Y(fft_d2[10]) );
  BUFX12 U463 ( .A(n3282), .Y(fft_d2[8]) );
  BUFX12 U464 ( .A(n3284), .Y(fft_d2[6]) );
  BUFX12 U465 ( .A(n3286), .Y(fft_d2[4]) );
  BUFX12 U466 ( .A(n3288), .Y(fft_d2[2]) );
  BUFX12 U467 ( .A(n3519), .Y(fft_d10[27]) );
  BUFX12 U468 ( .A(n3521), .Y(fft_d10[25]) );
  BUFX12 U469 ( .A(n3523), .Y(fft_d10[23]) );
  BUFX12 U470 ( .A(n3525), .Y(fft_d10[21]) );
  BUFX12 U471 ( .A(n3527), .Y(fft_d10[19]) );
  BUFX12 U472 ( .A(n3529), .Y(fft_d10[17]) );
  BUFX12 U473 ( .A(n3659), .Y(fft_d14[15]) );
  BUFX12 U474 ( .A(n3661), .Y(fft_d14[13]) );
  BUFX12 U475 ( .A(n3663), .Y(fft_d14[11]) );
  BUFX12 U476 ( .A(n3665), .Y(fft_d14[9]) );
  BUFX12 U477 ( .A(n3667), .Y(fft_d14[7]) );
  BUFX12 U478 ( .A(n3669), .Y(fft_d14[5]) );
  BUFX12 U479 ( .A(n3671), .Y(fft_d14[3]) );
  BUFX12 U480 ( .A(n3673), .Y(fft_d14[1]) );
  BUFX12 U481 ( .A(n3389), .Y(fft_d6[29]) );
  BUFX12 U482 ( .A(n3391), .Y(fft_d6[27]) );
  BUFX12 U483 ( .A(n3393), .Y(fft_d6[25]) );
  BUFX12 U484 ( .A(n3395), .Y(fft_d6[23]) );
  BUFX12 U485 ( .A(n3397), .Y(fft_d6[21]) );
  BUFX12 U486 ( .A(n3399), .Y(fft_d6[19]) );
  BUFX12 U487 ( .A(n3401), .Y(fft_d6[17]) );
  BUFX12 U488 ( .A(n3531), .Y(fft_d10[15]) );
  BUFX12 U489 ( .A(n3533), .Y(fft_d10[13]) );
  BUFX12 U490 ( .A(n3535), .Y(fft_d10[11]) );
  BUFX12 U491 ( .A(n3537), .Y(fft_d10[9]) );
  BUFX12 U492 ( .A(n3539), .Y(fft_d10[7]) );
  BUFX12 U493 ( .A(n3541), .Y(fft_d10[5]) );
  BUFX12 U494 ( .A(n3543), .Y(fft_d10[3]) );
  BUFX12 U495 ( .A(n3545), .Y(fft_d10[1]) );
  BUFX12 U496 ( .A(n3261), .Y(fft_d2[29]) );
  BUFX12 U497 ( .A(n3263), .Y(fft_d2[27]) );
  BUFX12 U498 ( .A(n3265), .Y(fft_d2[25]) );
  BUFX12 U499 ( .A(n3267), .Y(fft_d2[23]) );
  BUFX12 U500 ( .A(n3269), .Y(fft_d2[21]) );
  BUFX12 U501 ( .A(n3271), .Y(fft_d2[19]) );
  BUFX12 U502 ( .A(n3273), .Y(fft_d2[17]) );
  BUFX12 U503 ( .A(n3275), .Y(fft_d2[15]) );
  BUFX12 U504 ( .A(n3405), .Y(fft_d6[13]) );
  BUFX12 U505 ( .A(n3407), .Y(fft_d6[11]) );
  BUFX12 U506 ( .A(n3409), .Y(fft_d6[9]) );
  BUFX12 U507 ( .A(n3411), .Y(fft_d6[7]) );
  BUFX12 U508 ( .A(n3413), .Y(fft_d6[5]) );
  BUFX12 U509 ( .A(n3415), .Y(fft_d6[3]) );
  BUFX12 U510 ( .A(n3417), .Y(fft_d6[1]) );
  BUFX12 U511 ( .A(n3518), .Y(fft_d10[28]) );
  BUFX12 U512 ( .A(n3520), .Y(fft_d10[26]) );
  BUFX12 U513 ( .A(n3522), .Y(fft_d10[24]) );
  BUFX12 U514 ( .A(n3524), .Y(fft_d10[22]) );
  BUFX12 U515 ( .A(n3526), .Y(fft_d10[20]) );
  BUFX12 U516 ( .A(n3528), .Y(fft_d10[18]) );
  BUFX12 U517 ( .A(n3530), .Y(fft_d10[16]) );
  BUFX12 U518 ( .A(n3660), .Y(fft_d14[14]) );
  BUFX12 U519 ( .A(n3662), .Y(fft_d14[12]) );
  BUFX12 U520 ( .A(n3664), .Y(fft_d14[10]) );
  BUFX12 U521 ( .A(n3666), .Y(fft_d14[8]) );
  BUFX12 U522 ( .A(n3668), .Y(fft_d14[6]) );
  BUFX12 U523 ( .A(n3670), .Y(fft_d14[4]) );
  BUFX12 U524 ( .A(n3672), .Y(fft_d14[2]) );
  BUFX12 U525 ( .A(n3674), .Y(fft_d14[0]) );
  BUFX12 U526 ( .A(n3418), .Y(fft_d6[0]) );
  BUFX20 U527 ( .A(n3730), .Y(fft_d0[0]) );
  BUFX12 U528 ( .A(n3228), .Y(fft_d1[30]) );
  BUFX12 U529 ( .A(n3485), .Y(fft_d9[29]) );
  BUFX12 U530 ( .A(n3358), .Y(fft_d5[28]) );
  BUFX12 U531 ( .A(n3360), .Y(fft_d5[26]) );
  BUFX12 U532 ( .A(n3362), .Y(fft_d5[24]) );
  BUFX12 U533 ( .A(n3364), .Y(fft_d5[22]) );
  BUFX12 U534 ( .A(n3366), .Y(fft_d5[20]) );
  BUFX12 U535 ( .A(n3368), .Y(fft_d5[18]) );
  BUFX12 U536 ( .A(n3370), .Y(fft_d5[16]) );
  BUFX12 U537 ( .A(n3500), .Y(fft_d9[14]) );
  BUFX12 U538 ( .A(n3502), .Y(fft_d9[12]) );
  BUFX12 U539 ( .A(n3504), .Y(fft_d9[10]) );
  BUFX12 U540 ( .A(n3506), .Y(fft_d9[8]) );
  BUFX12 U541 ( .A(n3508), .Y(fft_d9[6]) );
  BUFX12 U542 ( .A(n3510), .Y(fft_d9[4]) );
  BUFX12 U543 ( .A(n3512), .Y(fft_d9[2]) );
  BUFX12 U544 ( .A(n3514), .Y(fft_d9[0]) );
  BUFX16 U545 ( .A(n3710), .Y(fft_d0[28]) );
  BUFX16 U546 ( .A(n3722), .Y(fft_d0[12]) );
  BUFX16 U547 ( .A(n3712), .Y(fft_d0[26]) );
  BUFX16 U548 ( .A(n3724), .Y(fft_d0[10]) );
  BUFX12 U549 ( .A(n3646), .Y(fft_d14[28]) );
  BUFX12 U550 ( .A(n3648), .Y(fft_d14[26]) );
  BUFX12 U551 ( .A(n3650), .Y(fft_d14[24]) );
  BUFX12 U552 ( .A(n3652), .Y(fft_d14[22]) );
  BUFX12 U553 ( .A(n3654), .Y(fft_d14[20]) );
  BUFX12 U554 ( .A(n3656), .Y(fft_d14[18]) );
  BUFX12 U555 ( .A(n3658), .Y(fft_d14[16]) );
  BUFX12 U556 ( .A(n3403), .Y(fft_d6[15]) );
  BUFX12 U557 ( .A(n3277), .Y(fft_d2[13]) );
  BUFX12 U558 ( .A(n3279), .Y(fft_d2[11]) );
  BUFX12 U559 ( .A(n3281), .Y(fft_d2[9]) );
  BUFX12 U560 ( .A(n3283), .Y(fft_d2[7]) );
  BUFX12 U561 ( .A(n3285), .Y(fft_d2[5]) );
  BUFX12 U562 ( .A(n3287), .Y(fft_d2[3]) );
  BUFX12 U563 ( .A(n3289), .Y(fft_d2[1]) );
  BUFX12 U564 ( .A(n3611), .Y(fft_d13[31]) );
  BUFX12 U565 ( .A(n3483), .Y(fft_d9[31]) );
  BUFX12 U566 ( .A(n3355), .Y(fft_d5[31]) );
  BUFX12 U567 ( .A(n3227), .Y(fft_d1[31]) );
  BUFX12 U568 ( .A(n3612), .Y(fft_d13[30]) );
  BUFX12 U569 ( .A(n3484), .Y(fft_d9[30]) );
  BUFX12 U570 ( .A(n3356), .Y(fft_d5[30]) );
  BUFX12 U571 ( .A(n3613), .Y(fft_d13[29]) );
  BUFX12 U572 ( .A(n3453), .Y(fft_d8[29]) );
  BUFX12 U573 ( .A(n3325), .Y(fft_d4[29]) );
  BUFX12 U574 ( .A(n3582), .Y(fft_d12[28]) );
  BUFX12 U575 ( .A(n3486), .Y(fft_d9[28]) );
  BUFX12 U576 ( .A(n3326), .Y(fft_d4[28]) );
  BUFX12 U577 ( .A(n3583), .Y(fft_d12[27]) );
  BUFX12 U578 ( .A(n3455), .Y(fft_d8[27]) );
  BUFX12 U579 ( .A(n3327), .Y(fft_d4[27]) );
  BUFX12 U580 ( .A(n3584), .Y(fft_d12[26]) );
  BUFX12 U581 ( .A(n3488), .Y(fft_d9[26]) );
  BUFX12 U582 ( .A(n3328), .Y(fft_d4[26]) );
  BUFX12 U583 ( .A(n3585), .Y(fft_d12[25]) );
  BUFX12 U584 ( .A(n3457), .Y(fft_d8[25]) );
  BUFX12 U585 ( .A(n3329), .Y(fft_d4[25]) );
  BUFX12 U586 ( .A(n3586), .Y(fft_d12[24]) );
  BUFX12 U587 ( .A(n3490), .Y(fft_d9[24]) );
  BUFX12 U588 ( .A(n3330), .Y(fft_d4[24]) );
  BUFX12 U589 ( .A(n3587), .Y(fft_d12[23]) );
  BUFX12 U590 ( .A(n3459), .Y(fft_d8[23]) );
  BUFX12 U591 ( .A(n3331), .Y(fft_d4[23]) );
  BUFX12 U592 ( .A(n3588), .Y(fft_d12[22]) );
  BUFX12 U593 ( .A(n3492), .Y(fft_d9[22]) );
  BUFX12 U594 ( .A(n3332), .Y(fft_d4[22]) );
  BUFX12 U595 ( .A(n3589), .Y(fft_d12[21]) );
  BUFX12 U596 ( .A(n3461), .Y(fft_d8[21]) );
  BUFX12 U597 ( .A(n3333), .Y(fft_d4[21]) );
  BUFX12 U598 ( .A(n3590), .Y(fft_d12[20]) );
  BUFX12 U599 ( .A(n3494), .Y(fft_d9[20]) );
  BUFX12 U600 ( .A(n3334), .Y(fft_d4[20]) );
  BUFX12 U601 ( .A(n3591), .Y(fft_d12[19]) );
  BUFX12 U602 ( .A(n3463), .Y(fft_d8[19]) );
  BUFX12 U603 ( .A(n3335), .Y(fft_d4[19]) );
  BUFX12 U604 ( .A(n3592), .Y(fft_d12[18]) );
  BUFX12 U605 ( .A(n3496), .Y(fft_d9[18]) );
  BUFX12 U606 ( .A(n3336), .Y(fft_d4[18]) );
  BUFX12 U607 ( .A(n3593), .Y(fft_d12[17]) );
  BUFX12 U608 ( .A(n3465), .Y(fft_d8[17]) );
  BUFX12 U609 ( .A(n3337), .Y(fft_d4[17]) );
  BUFX12 U610 ( .A(n3594), .Y(fft_d12[16]) );
  BUFX12 U611 ( .A(n3498), .Y(fft_d9[16]) );
  BUFX12 U612 ( .A(n3338), .Y(fft_d4[16]) );
  BUFX12 U613 ( .A(n3595), .Y(fft_d12[15]) );
  BUFX12 U614 ( .A(n3467), .Y(fft_d8[15]) );
  BUFX12 U615 ( .A(n3339), .Y(fft_d4[15]) );
  BUFX12 U616 ( .A(n3243), .Y(fft_d1[15]) );
  BUFX12 U617 ( .A(n3628), .Y(fft_d13[14]) );
  BUFX12 U618 ( .A(n3468), .Y(fft_d8[14]) );
  BUFX12 U619 ( .A(n3340), .Y(fft_d4[14]) );
  BUFX12 U620 ( .A(n3597), .Y(fft_d12[13]) );
  BUFX12 U621 ( .A(n3469), .Y(fft_d8[13]) );
  BUFX12 U622 ( .A(n3341), .Y(fft_d4[13]) );
  BUFX12 U623 ( .A(n3630), .Y(fft_d13[12]) );
  BUFX12 U624 ( .A(n3470), .Y(fft_d8[12]) );
  BUFX12 U625 ( .A(n3342), .Y(fft_d4[12]) );
  BUFX12 U626 ( .A(n3599), .Y(fft_d12[11]) );
  BUFX12 U627 ( .A(n3471), .Y(fft_d8[11]) );
  BUFX12 U628 ( .A(n3343), .Y(fft_d4[11]) );
  BUFX12 U629 ( .A(n3632), .Y(fft_d13[10]) );
  BUFX12 U630 ( .A(n3472), .Y(fft_d8[10]) );
  BUFX12 U631 ( .A(n3344), .Y(fft_d4[10]) );
  BUFX12 U632 ( .A(n3601), .Y(fft_d12[9]) );
  BUFX12 U633 ( .A(n3473), .Y(fft_d8[9]) );
  BUFX12 U634 ( .A(n3345), .Y(fft_d4[9]) );
  BUFX12 U635 ( .A(n3634), .Y(fft_d13[8]) );
  BUFX12 U636 ( .A(n3474), .Y(fft_d8[8]) );
  BUFX12 U637 ( .A(n3346), .Y(fft_d4[8]) );
  BUFX12 U638 ( .A(n3603), .Y(fft_d12[7]) );
  BUFX12 U639 ( .A(n3475), .Y(fft_d8[7]) );
  BUFX12 U640 ( .A(n3347), .Y(fft_d4[7]) );
  BUFX12 U641 ( .A(n3636), .Y(fft_d13[6]) );
  BUFX12 U642 ( .A(n3476), .Y(fft_d8[6]) );
  BUFX12 U643 ( .A(n3348), .Y(fft_d4[6]) );
  BUFX12 U644 ( .A(n3605), .Y(fft_d12[5]) );
  BUFX12 U645 ( .A(n3477), .Y(fft_d8[5]) );
  BUFX12 U646 ( .A(n3349), .Y(fft_d4[5]) );
  BUFX12 U647 ( .A(n3638), .Y(fft_d13[4]) );
  BUFX12 U648 ( .A(n3478), .Y(fft_d8[4]) );
  BUFX12 U649 ( .A(n3350), .Y(fft_d4[4]) );
  BUFX12 U650 ( .A(n3607), .Y(fft_d12[3]) );
  BUFX12 U651 ( .A(n3479), .Y(fft_d8[3]) );
  BUFX12 U652 ( .A(n3351), .Y(fft_d4[3]) );
  BUFX12 U653 ( .A(n3640), .Y(fft_d13[2]) );
  BUFX12 U654 ( .A(n3480), .Y(fft_d8[2]) );
  BUFX12 U655 ( .A(n3352), .Y(fft_d4[2]) );
  BUFX12 U656 ( .A(n3609), .Y(fft_d12[1]) );
  BUFX12 U657 ( .A(n3481), .Y(fft_d8[1]) );
  BUFX12 U658 ( .A(n3353), .Y(fft_d4[1]) );
  BUFX12 U659 ( .A(n3642), .Y(fft_d13[0]) );
  BUFX12 U660 ( .A(n3482), .Y(fft_d8[0]) );
  BUFX12 U661 ( .A(n3386), .Y(fft_d5[0]) );
  BUFX12 U662 ( .A(n3258), .Y(fft_d1[0]) );
  BUFX12 U663 ( .A(n3547), .Y(fft_d11[31]) );
  BUFX12 U664 ( .A(n3419), .Y(fft_d7[31]) );
  BUFX12 U665 ( .A(n3291), .Y(fft_d3[31]) );
  BUFX12 U666 ( .A(n3676), .Y(fft_d15[30]) );
  BUFX12 U667 ( .A(n3548), .Y(fft_d11[30]) );
  BUFX12 U668 ( .A(n3420), .Y(fft_d7[30]) );
  BUFX12 U669 ( .A(n3292), .Y(fft_d3[30]) );
  BUFX12 U670 ( .A(n3677), .Y(fft_d15[29]) );
  BUFX12 U671 ( .A(n3549), .Y(fft_d11[29]) );
  BUFX12 U672 ( .A(n3422), .Y(fft_d7[28]) );
  BUFX12 U673 ( .A(n3424), .Y(fft_d7[26]) );
  BUFX12 U674 ( .A(n3426), .Y(fft_d7[24]) );
  BUFX12 U675 ( .A(n3428), .Y(fft_d7[22]) );
  BUFX12 U676 ( .A(n3430), .Y(fft_d7[20]) );
  BUFX12 U677 ( .A(n3432), .Y(fft_d7[18]) );
  BUFX12 U678 ( .A(n3434), .Y(fft_d7[16]) );
  BUFX12 U679 ( .A(n3564), .Y(fft_d11[14]) );
  BUFX12 U680 ( .A(n3566), .Y(fft_d11[12]) );
  BUFX12 U681 ( .A(n3568), .Y(fft_d11[10]) );
  BUFX12 U682 ( .A(n3570), .Y(fft_d11[8]) );
  BUFX12 U683 ( .A(n3572), .Y(fft_d11[6]) );
  BUFX12 U684 ( .A(n3574), .Y(fft_d11[4]) );
  BUFX12 U685 ( .A(n3576), .Y(fft_d11[2]) );
  BUFX12 U686 ( .A(n3578), .Y(fft_d11[0]) );
  BUFX12 U687 ( .A(n3322), .Y(fft_d3[0]) );
  BUFX16 U688 ( .A(n3708), .Y(fft_d0[30]) );
  BUFX16 U689 ( .A(n3720), .Y(fft_d0[14]) );
  BUFX16 U690 ( .A(n3711), .Y(fft_d0[27]) );
  BUFX16 U691 ( .A(n3709), .Y(fft_d0[29]) );
  BUFX16 U692 ( .A(n3721), .Y(fft_d0[13]) );
  BUFX12 U693 ( .A(n3579), .Y(fft_d12[31]) );
  BUFX12 U694 ( .A(n3451), .Y(fft_d8[31]) );
  BUFX12 U695 ( .A(n3323), .Y(fft_d4[31]) );
  BUFX12 U696 ( .A(n3580), .Y(fft_d12[30]) );
  BUFX12 U697 ( .A(n3452), .Y(fft_d8[30]) );
  BUFX12 U698 ( .A(n3324), .Y(fft_d4[30]) );
  BUFX12 U699 ( .A(n3581), .Y(fft_d12[29]) );
  BUFX12 U700 ( .A(n3357), .Y(fft_d5[29]) );
  BUFX12 U701 ( .A(n3229), .Y(fft_d1[29]) );
  BUFX12 U702 ( .A(n3614), .Y(fft_d13[28]) );
  BUFX12 U703 ( .A(n3454), .Y(fft_d8[28]) );
  BUFX12 U704 ( .A(n3230), .Y(fft_d1[28]) );
  BUFX12 U705 ( .A(n3615), .Y(fft_d13[27]) );
  BUFX12 U706 ( .A(n3487), .Y(fft_d9[27]) );
  BUFX12 U707 ( .A(n3359), .Y(fft_d5[27]) );
  BUFX12 U708 ( .A(n3231), .Y(fft_d1[27]) );
  BUFX12 U709 ( .A(n3616), .Y(fft_d13[26]) );
  BUFX12 U710 ( .A(n3456), .Y(fft_d8[26]) );
  BUFX12 U711 ( .A(n3232), .Y(fft_d1[26]) );
  BUFX12 U712 ( .A(n3617), .Y(fft_d13[25]) );
  BUFX12 U713 ( .A(n3489), .Y(fft_d9[25]) );
  BUFX12 U714 ( .A(n3361), .Y(fft_d5[25]) );
  BUFX12 U715 ( .A(n3233), .Y(fft_d1[25]) );
  BUFX12 U716 ( .A(n3618), .Y(fft_d13[24]) );
  BUFX12 U717 ( .A(n3458), .Y(fft_d8[24]) );
  BUFX12 U718 ( .A(n3234), .Y(fft_d1[24]) );
  BUFX12 U719 ( .A(n3619), .Y(fft_d13[23]) );
  BUFX12 U720 ( .A(n3491), .Y(fft_d9[23]) );
  BUFX12 U721 ( .A(n3363), .Y(fft_d5[23]) );
  BUFX12 U722 ( .A(n3235), .Y(fft_d1[23]) );
  BUFX12 U723 ( .A(n3620), .Y(fft_d13[22]) );
  BUFX12 U724 ( .A(n3460), .Y(fft_d8[22]) );
  BUFX12 U725 ( .A(n3621), .Y(fft_d13[21]) );
  BUFX12 U726 ( .A(n3493), .Y(fft_d9[21]) );
  BUFX12 U727 ( .A(n3365), .Y(fft_d5[21]) );
  BUFX12 U728 ( .A(n3622), .Y(fft_d13[20]) );
  BUFX12 U729 ( .A(n3462), .Y(fft_d8[20]) );
  BUFX12 U730 ( .A(n3623), .Y(fft_d13[19]) );
  BUFX12 U731 ( .A(n3495), .Y(fft_d9[19]) );
  BUFX12 U732 ( .A(n3367), .Y(fft_d5[19]) );
  BUFX12 U733 ( .A(n3624), .Y(fft_d13[18]) );
  BUFX12 U734 ( .A(n3464), .Y(fft_d8[18]) );
  BUFX12 U735 ( .A(n3240), .Y(fft_d1[18]) );
  BUFX12 U736 ( .A(n3625), .Y(fft_d13[17]) );
  BUFX12 U737 ( .A(n3497), .Y(fft_d9[17]) );
  BUFX12 U738 ( .A(n3369), .Y(fft_d5[17]) );
  BUFX12 U739 ( .A(n3626), .Y(fft_d13[16]) );
  BUFX12 U740 ( .A(n3466), .Y(fft_d8[16]) );
  BUFX12 U741 ( .A(n3242), .Y(fft_d1[16]) );
  BUFX12 U742 ( .A(n3627), .Y(fft_d13[15]) );
  BUFX12 U743 ( .A(n3499), .Y(fft_d9[15]) );
  BUFX12 U744 ( .A(n3371), .Y(fft_d5[15]) );
  BUFX12 U745 ( .A(n3596), .Y(fft_d12[14]) );
  BUFX12 U746 ( .A(n3372), .Y(fft_d5[14]) );
  BUFX12 U747 ( .A(n3244), .Y(fft_d1[14]) );
  BUFX12 U748 ( .A(n3629), .Y(fft_d13[13]) );
  BUFX12 U749 ( .A(n3501), .Y(fft_d9[13]) );
  BUFX12 U750 ( .A(n3373), .Y(fft_d5[13]) );
  BUFX12 U751 ( .A(n3245), .Y(fft_d1[13]) );
  BUFX12 U752 ( .A(n3598), .Y(fft_d12[12]) );
  BUFX12 U753 ( .A(n3374), .Y(fft_d5[12]) );
  BUFX12 U754 ( .A(n3246), .Y(fft_d1[12]) );
  BUFX12 U755 ( .A(n3631), .Y(fft_d13[11]) );
  BUFX12 U756 ( .A(n3503), .Y(fft_d9[11]) );
  BUFX12 U757 ( .A(n3375), .Y(fft_d5[11]) );
  BUFX12 U758 ( .A(n3247), .Y(fft_d1[11]) );
  BUFX12 U759 ( .A(n3600), .Y(fft_d12[10]) );
  BUFX12 U760 ( .A(n3376), .Y(fft_d5[10]) );
  BUFX12 U761 ( .A(n3248), .Y(fft_d1[10]) );
  BUFX12 U762 ( .A(n3633), .Y(fft_d13[9]) );
  BUFX12 U763 ( .A(n3505), .Y(fft_d9[9]) );
  BUFX12 U764 ( .A(n3377), .Y(fft_d5[9]) );
  BUFX12 U765 ( .A(n3249), .Y(fft_d1[9]) );
  BUFX12 U766 ( .A(n3602), .Y(fft_d12[8]) );
  BUFX12 U767 ( .A(n3378), .Y(fft_d5[8]) );
  BUFX12 U768 ( .A(n3250), .Y(fft_d1[8]) );
  BUFX12 U769 ( .A(n3635), .Y(fft_d13[7]) );
  BUFX12 U770 ( .A(n3507), .Y(fft_d9[7]) );
  BUFX12 U771 ( .A(n3379), .Y(fft_d5[7]) );
  BUFX12 U772 ( .A(n3251), .Y(fft_d1[7]) );
  BUFX12 U773 ( .A(n3604), .Y(fft_d12[6]) );
  BUFX12 U774 ( .A(n3380), .Y(fft_d5[6]) );
  BUFX12 U775 ( .A(n3637), .Y(fft_d13[5]) );
  BUFX12 U776 ( .A(n3509), .Y(fft_d9[5]) );
  BUFX12 U777 ( .A(n3381), .Y(fft_d5[5]) );
  BUFX12 U778 ( .A(n3606), .Y(fft_d12[4]) );
  BUFX12 U779 ( .A(n3382), .Y(fft_d5[4]) );
  BUFX12 U780 ( .A(n3639), .Y(fft_d13[3]) );
  BUFX12 U781 ( .A(n3511), .Y(fft_d9[3]) );
  BUFX12 U782 ( .A(n3383), .Y(fft_d5[3]) );
  BUFX12 U783 ( .A(n3608), .Y(fft_d12[2]) );
  BUFX12 U784 ( .A(n3384), .Y(fft_d5[2]) );
  BUFX12 U785 ( .A(n3256), .Y(fft_d1[2]) );
  BUFX12 U786 ( .A(n3641), .Y(fft_d13[1]) );
  BUFX12 U787 ( .A(n3513), .Y(fft_d9[1]) );
  BUFX12 U788 ( .A(n3385), .Y(fft_d5[1]) );
  BUFX12 U789 ( .A(n3610), .Y(fft_d12[0]) );
  BUFX12 U790 ( .A(n3354), .Y(fft_d4[0]) );
  BUFX12 U791 ( .A(n3239), .Y(fft_d1[19]) );
  BUFX12 U792 ( .A(n3241), .Y(fft_d1[17]) );
  BUFX12 U793 ( .A(n3257), .Y(fft_d1[1]) );
  BUFX12 U794 ( .A(n3255), .Y(fft_d1[3]) );
  BUFX12 U795 ( .A(n3238), .Y(fft_d1[20]) );
  BUFX12 U796 ( .A(n3254), .Y(fft_d1[4]) );
  BUFX12 U797 ( .A(n3237), .Y(fft_d1[21]) );
  BUFX12 U798 ( .A(n3253), .Y(fft_d1[5]) );
  BUFX12 U799 ( .A(n3236), .Y(fft_d1[22]) );
  BUFX12 U800 ( .A(n3252), .Y(fft_d1[6]) );
  BUFX12 U801 ( .A(n3515), .Y(fft_d10[31]) );
  BUFX12 U802 ( .A(n3387), .Y(fft_d6[31]) );
  BUFX12 U803 ( .A(n3259), .Y(fft_d2[31]) );
  BUFX12 U804 ( .A(n3644), .Y(fft_d14[30]) );
  BUFX12 U805 ( .A(n3516), .Y(fft_d10[30]) );
  BUFX12 U806 ( .A(n3388), .Y(fft_d6[30]) );
  BUFX12 U807 ( .A(n3260), .Y(fft_d2[30]) );
  BUFX12 U808 ( .A(n3645), .Y(fft_d14[29]) );
  BUFX12 U809 ( .A(n3517), .Y(fft_d10[29]) );
  BUFX12 U810 ( .A(n3390), .Y(fft_d6[28]) );
  BUFX12 U811 ( .A(n3392), .Y(fft_d6[26]) );
  BUFX12 U812 ( .A(n3394), .Y(fft_d6[24]) );
  BUFX12 U813 ( .A(n3396), .Y(fft_d6[22]) );
  BUFX12 U814 ( .A(n3398), .Y(fft_d6[20]) );
  BUFX12 U815 ( .A(n3400), .Y(fft_d6[18]) );
  BUFX12 U816 ( .A(n3402), .Y(fft_d6[16]) );
  BUFX12 U817 ( .A(n3532), .Y(fft_d10[14]) );
  BUFX12 U818 ( .A(n3534), .Y(fft_d10[12]) );
  BUFX12 U819 ( .A(n3536), .Y(fft_d10[10]) );
  BUFX12 U820 ( .A(n3538), .Y(fft_d10[8]) );
  BUFX12 U821 ( .A(n3540), .Y(fft_d10[6]) );
  BUFX12 U822 ( .A(n3542), .Y(fft_d10[4]) );
  BUFX12 U823 ( .A(n3544), .Y(fft_d10[2]) );
  BUFX12 U824 ( .A(n3546), .Y(fft_d10[0]) );
  BUFX12 U825 ( .A(n3290), .Y(fft_d2[0]) );
  INVX12 U826 ( .A(n7160), .Y(fft_valid) );
  BUFX16 U827 ( .A(n3707), .Y(fft_d0[31]) );
  BUFX16 U828 ( .A(n3719), .Y(fft_d0[15]) );
  CLKINVX12 U829 ( .A(n3728), .Y(n7200) );
  CLKINVX20 U830 ( .A(n7200), .Y(fft_d0[6]) );
  CLKINVX12 U831 ( .A(n3716), .Y(n7220) );
  CLKINVX20 U832 ( .A(n7220), .Y(fft_d0[22]) );
  NAND3BX2 U833 ( .AN(n1790), .B(n109), .C(n177), .Y(n10500) );
  INVX3 U834 ( .A(mul_2_Wn[14]), .Y(n2863) );
  OA22XL U835 ( .A0(n19), .A1(n2943), .B0(n185), .B1(n2942), .Y(n2947) );
  CLKINVX1 U836 ( .A(stg_reg[113]), .Y(n2846) );
  OA22X1 U837 ( .A0(n906), .A1(n2939), .B0(n46), .B1(n2940), .Y(n2937) );
  OA22XL U838 ( .A0(n47), .A1(n3034), .B0(n9630), .B1(n3033), .Y(n3038) );
  CLKINVX1 U839 ( .A(stg_reg[97]), .Y(n3049) );
  OA22XL U840 ( .A0(n906), .A1(n2913), .B0(n49), .B1(n2914), .Y(n2911) );
  INVX3 U841 ( .A(n841), .Y(n3055) );
  NAND2X1 U842 ( .A(n7320), .B(n2861), .Y(mul_0_Wn[13]) );
  OA22X1 U843 ( .A0(n908), .A1(n2965), .B0(n20), .B1(n2966), .Y(n2963) );
  CLKINVX1 U844 ( .A(stg_reg[96]), .Y(n3063) );
  INVX1 U845 ( .A(stg_reg[4]), .Y(n3009) );
  INVX1 U846 ( .A(stg_reg[116]), .Y(n2816) );
  CLKINVX1 U847 ( .A(stg_reg[112]), .Y(n2856) );
  NAND2XL U848 ( .A(n195), .B(n7300), .Y(mul_0_Wn[11]) );
  CLKBUFX2 U849 ( .A(n903), .Y(n907) );
  CLKBUFX2 U850 ( .A(n3072), .Y(n9190) );
  OA22XL U851 ( .A0(n908), .A1(n2926), .B0(n50), .B1(n2927), .Y(n2924) );
  OA22XL U852 ( .A0(n906), .A1(n2900), .B0(n47), .B1(n2901), .Y(n2898) );
  OA22XL U853 ( .A0(n9280), .A1(n2762), .B0(n9220), .B1(n2761), .Y(n2769) );
  OA22XL U854 ( .A0(n46), .A1(n2764), .B0(n187), .B1(n2763), .Y(n2768) );
  OA22XL U855 ( .A0(n77), .A1(n2766), .B0(n10460), .B1(n2765), .Y(n2767) );
  CLKINVX1 U856 ( .A(stg_reg[16]), .Y(n2855) );
  INVX1 U857 ( .A(stg_reg[102]), .Y(n2984) );
  CLKINVX1 U858 ( .A(stg_reg[108]), .Y(n2906) );
  CLKINVX1 U859 ( .A(stg_reg[109]), .Y(n2893) );
  CLKINVX1 U860 ( .A(stg_reg[110]), .Y(n2881) );
  CLKINVX1 U861 ( .A(stg_reg[122]), .Y(n2756) );
  CLKINVX1 U862 ( .A(stg_reg[125]), .Y(n2726) );
  CLKINVX1 U863 ( .A(stg_reg[126]), .Y(n2716) );
  INVX1 U864 ( .A(stg_reg[26]), .Y(n2755) );
  INVX1 U865 ( .A(stg_reg[27]), .Y(n2745) );
  CLKINVX1 U866 ( .A(stg_reg[12]), .Y(n2905) );
  CLKINVX1 U867 ( .A(stg_reg[13]), .Y(n2892) );
  CLKINVX1 U868 ( .A(stg_reg[30]), .Y(n2715) );
  CLKINVX1 U869 ( .A(stg_reg[14]), .Y(n2880) );
  CLKBUFX3 U870 ( .A(n9820), .Y(n9760) );
  NAND2X2 U871 ( .A(n7320), .B(n9680), .Y(mul_0_Wn[15]) );
  OA22X1 U872 ( .A0(n47), .A1(n2398), .B0(n191), .B1(n2889), .Y(n2397) );
  AOI2BB1X1 U873 ( .A0N(n852), .A1N(n2573), .B0(n832), .Y(n2570) );
  AOI2BB1X1 U874 ( .A0N(n851), .A1N(n2582), .B0(n833), .Y(n2579) );
  AOI2BB1X1 U875 ( .A0N(n851), .A1N(n2591), .B0(n834), .Y(n2588) );
  AOI2BB1X1 U876 ( .A0N(n851), .A1N(n2600), .B0(n823), .Y(n2597) );
  OA22XL U877 ( .A0(n49), .A1(n2969), .B0(n203), .B1(n2968), .Y(n2973) );
  OA22XL U878 ( .A0(n48), .A1(n3021), .B0(n185), .B1(n3020), .Y(n3025) );
  AOI2BB1X1 U879 ( .A0N(n851), .A1N(n2609), .B0(n824), .Y(n2606) );
  AOI2BB1X1 U880 ( .A0N(n851), .A1N(n2618), .B0(n825), .Y(n2615) );
  AOI2BB1X1 U881 ( .A0N(n851), .A1N(n2627), .B0(n826), .Y(n2624) );
  OAI221X1 U882 ( .A0(n9790), .A1(n2854), .B0(n46), .B1(n2853), .C0(n2386), 
        .Y(stg2_real_Wn[32]) );
  NAND2XL U883 ( .A(n10530), .B(n10360), .Y(n7270) );
  AOI222XL U884 ( .A0(stg_reg[40]), .A1(n861), .B0(n914), .B1(stg_reg[72]), 
        .C0(n905), .C1(n1576), .Y(n2962) );
  INVX1 U885 ( .A(stg_reg[104]), .Y(n2958) );
  INVX1 U886 ( .A(stg_reg[120]), .Y(n2776) );
  INVX1 U887 ( .A(stg_reg[100]), .Y(n3010) );
  INVX1 U888 ( .A(stg_reg[6]), .Y(n2983) );
  INVXL U889 ( .A(stg_reg[77]), .Y(n3088) );
  INVXL U890 ( .A(stg_reg[93]), .Y(n1306) );
  CLKINVX3 U891 ( .A(mul_o_sub[19]), .Y(n2663) );
  CLKBUFX2 U892 ( .A(n9820), .Y(n9780) );
  CLKBUFX2 U893 ( .A(n9790), .Y(n9770) );
  NAND2X4 U894 ( .A(n7300), .B(n10540), .Y(mul_2_Wn_11) );
  CLKBUFX2 U895 ( .A(n3148), .Y(n9820) );
  CLKBUFX2 U896 ( .A(n3148), .Y(n9810) );
  AND2XL U897 ( .A(n1287), .B(n10540), .Y(n7310) );
  CLKBUFX2 U898 ( .A(n7260), .Y(n916) );
  INVX1 U899 ( .A(stg4_img[30]), .Y(n2879) );
  INVX1 U900 ( .A(stg4_img[14]), .Y(n2472) );
  INVX1 U901 ( .A(stg4_img[31]), .Y(n3083) );
  NAND3BXL U902 ( .AN(n1420), .B(n2864), .C(n909), .Y(n10590) );
  NAND3BXL U903 ( .AN(mul_0_Wn[13]), .B(n1417), .C(n866), .Y(n1285) );
  NAND3BXL U904 ( .AN(n1420), .B(n7320), .C(n9200), .Y(n1421) );
  NAND3BXL U905 ( .AN(mul_2_Wn_11), .B(n1417), .C(n917), .Y(n1418) );
  CLKBUFX2 U906 ( .A(n867), .Y(n866) );
  CLKBUFX2 U907 ( .A(n867), .Y(n865) );
  CLKBUFX2 U908 ( .A(n866), .Y(n864) );
  NAND2XL U909 ( .A(n10460), .B(n7320), .Y(mul_0_Wn[12]) );
  CLKBUFX2 U910 ( .A(n9210), .Y(n9200) );
  INVX1 U911 ( .A(stg4_real[31]), .Y(n3070) );
  NAND3BXL U912 ( .AN(n1284), .B(n7300), .C(n9340), .Y(n1420) );
  NAND3BXL U913 ( .AN(n1284), .B(n1301), .C(n9280), .Y(n10580) );
  CLKBUFX2 U914 ( .A(n906), .Y(n908) );
  XNOR2X1 U915 ( .A(stg2_img_11__15_), .B(n7480), .Y(stg2_img_15__15_) );
  XNOR2X1 U916 ( .A(stg2_img_10__15_), .B(n7890), .Y(stg2_img_14__15_) );
  XNOR2X1 U917 ( .A(stg2_img_9__15_), .B(n7900), .Y(stg2_img_13__15_) );
  OA22XL U918 ( .A0(n50), .A1(n2402), .B0(n195), .B1(n2900), .Y(n2401) );
  OA22XL U919 ( .A0(n9200), .A1(n2900), .B0(n51), .B1(n2482), .Y(n2481) );
  AOI2BB2XL U920 ( .B0(stg2_img_15__13_), .B1(n872), .A0N(n2889), .A1N(n851), 
        .Y(n2475) );
  AOI2BB2XL U921 ( .B0(stg2_img_15__12_), .B1(n872), .A0N(n2900), .A1N(n851), 
        .Y(n2480) );
  OA22XL U922 ( .A0(n47), .A1(n3047), .B0(n199), .B1(n3046), .Y(n3051) );
  OA22XL U923 ( .A0(n50), .A1(n2995), .B0(n9630), .B1(n2994), .Y(n2999) );
  OA22XL U924 ( .A0(n9280), .A1(n2822), .B0(n3072), .B1(n2821), .Y(n2829) );
  OA22XL U925 ( .A0(n9280), .A1(n2842), .B0(n3072), .B1(n2841), .Y(n2849) );
  OA22XL U926 ( .A0(n9280), .A1(n2802), .B0(n3072), .B1(n2801), .Y(n2809) );
  OA22XL U927 ( .A0(n9280), .A1(n2782), .B0(n3072), .B1(n2781), .Y(n2789) );
  OA22XL U928 ( .A0(n9280), .A1(n2832), .B0(n3072), .B1(n2831), .Y(n2839) );
  OA22XL U929 ( .A0(n9280), .A1(n2812), .B0(n9220), .B1(n2811), .Y(n2819) );
  OA22XL U930 ( .A0(n9280), .A1(n2792), .B0(n9210), .B1(n2791), .Y(n2799) );
  OA22XL U931 ( .A0(n9280), .A1(n2772), .B0(n9190), .B1(n2771), .Y(n2779) );
  OA22XL U932 ( .A0(n48), .A1(n2982), .B0(n207), .B1(n2981), .Y(n2986) );
  OA22XL U933 ( .A0(n52), .A1(n3008), .B0(n195), .B1(n3007), .Y(n3012) );
  OA22XL U934 ( .A0(n51), .A1(n2956), .B0(n197), .B1(n2955), .Y(n2960) );
  OA22XL U935 ( .A0(n20), .A1(n2904), .B0(n181), .B1(n2903), .Y(n2908) );
  OA22XL U936 ( .A0(n52), .A1(n2930), .B0(n195), .B1(n2929), .Y(n2934) );
  OA22XL U937 ( .A0(n51), .A1(n2406), .B0(n191), .B1(n2913), .Y(n2405) );
  OA22XL U938 ( .A0(n917), .A1(n2913), .B0(n51), .B1(n2487), .Y(n2486) );
  OA22XL U939 ( .A0(n20), .A1(n2410), .B0(n181), .B1(n2926), .Y(n2409) );
  OA22XL U940 ( .A0(n9200), .A1(n2926), .B0(n52), .B1(n2492), .Y(n2491) );
  OA22XL U941 ( .A0(n49), .A1(n2414), .B0(n193), .B1(n2939), .Y(n2413) );
  OA22XL U942 ( .A0(n917), .A1(n2939), .B0(n49), .B1(n2497), .Y(n2496) );
  OA22XL U943 ( .A0(n52), .A1(n2418), .B0(n195), .B1(n2952), .Y(n2417) );
  OA22XL U944 ( .A0(n906), .A1(n2952), .B0(n46), .B1(n2953), .Y(n2950) );
  OA22XL U945 ( .A0(n9190), .A1(n2952), .B0(n50), .B1(n2502), .Y(n2501) );
  AOI2BB2XL U946 ( .B0(stg2_img_15__11_), .B1(n872), .A0N(n2913), .A1N(n2687), 
        .Y(n2485) );
  AOI2BB2XL U947 ( .B0(stg2_img_15__10_), .B1(n872), .A0N(n2926), .A1N(n852), 
        .Y(n2490) );
  AOI2BB2XL U948 ( .B0(stg2_img_15__9_), .B1(n872), .A0N(n2939), .A1N(n851), 
        .Y(n2495) );
  AOI2BB2XL U949 ( .B0(stg2_img_15__8_), .B1(n872), .A0N(n2952), .A1N(n851), 
        .Y(n2500) );
  OA22XL U950 ( .A0(n9280), .A1(n2742), .B0(n3072), .B1(n2741), .Y(n2749) );
  OA22XL U951 ( .A0(n9280), .A1(n2852), .B0(n3072), .B1(n2851), .Y(n2859) );
  OA22XL U952 ( .A0(n9280), .A1(n2722), .B0(n3072), .B1(n2721), .Y(n2729) );
  OA22XL U953 ( .A0(n9280), .A1(n2713), .B0(n9220), .B1(n2712), .Y(n2719) );
  OA22XL U954 ( .A0(n94), .A1(n9280), .B0(n9200), .B1(n112), .Y(n2884) );
  OA22XL U955 ( .A0(n3098), .A1(n9280), .B0(n918), .B1(n2915), .Y(n2922) );
  OA22XL U956 ( .A0(n3147), .A1(n9280), .B0(n9210), .B1(n3059), .Y(n3066) );
  OA22XL U957 ( .A0(n3090), .A1(n9280), .B0(n9190), .B1(n108), .Y(n2896) );
  OA22XL U958 ( .A0(n9280), .A1(n2732), .B0(n3072), .B1(n2731), .Y(n2739) );
  OA22XL U959 ( .A0(n9280), .A1(n2752), .B0(n3072), .B1(n2751), .Y(n2759) );
  OAI221XL U960 ( .A0(n9760), .A1(n2832), .B0(n48), .B1(n115), .C0(n1400), .Y(
        stg2_real_Wn[18]) );
  OAI221XL U961 ( .A0(n9760), .A1(n2822), .B0(n46), .B1(n119), .C0(n1392), .Y(
        stg2_real_Wn[19]) );
  OAI221XL U962 ( .A0(n9760), .A1(n2842), .B0(n45), .B1(n116), .C0(n1408), .Y(
        stg2_real_Wn[17]) );
  OAI221XL U963 ( .A0(n9760), .A1(n2812), .B0(n20), .B1(n118), .C0(n1384), .Y(
        stg2_real_Wn[20]) );
  OAI221XL U964 ( .A0(n9780), .A1(n2844), .B0(n47), .B1(n2843), .C0(n2379), 
        .Y(stg2_real_Wn[33]) );
  OAI221XL U965 ( .A0(n9740), .A1(n2834), .B0(n51), .B1(n2833), .C0(n2372), 
        .Y(stg2_real_Wn[34]) );
  OAI221XL U966 ( .A0(n9770), .A1(n2824), .B0(n50), .B1(n2823), .C0(n2365), 
        .Y(stg2_real_Wn[35]) );
  OAI221XL U967 ( .A0(n9770), .A1(n2814), .B0(n48), .B1(n2813), .C0(n2358), 
        .Y(stg2_real_Wn[36]) );
  OA22XL U968 ( .A0(n205), .A1(n2816), .B0(n80), .B1(n2357), .Y(n2358) );
  OAI221XL U969 ( .A0(n9800), .A1(n2835), .B0(n46), .B1(n2831), .C0(n2677), 
        .Y(stg2_real_Wn[2]) );
  OAI221XL U970 ( .A0(n9750), .A1(n2825), .B0(n20), .B1(n2821), .C0(n2668), 
        .Y(stg2_real_Wn[3]) );
  OAI221XL U971 ( .A0(n9750), .A1(n2815), .B0(n52), .B1(n2811), .C0(n2659), 
        .Y(stg2_real_Wn[4]) );
  OAI221XL U972 ( .A0(n9750), .A1(n1274), .B0(n45), .B1(n1273), .C0(n1272), 
        .Y(stg2_real_Wn[49]) );
  OAI221XL U973 ( .A0(n9750), .A1(n1265), .B0(n52), .B1(n1264), .C0(n1263), 
        .Y(stg2_real_Wn[50]) );
  OAI221XL U974 ( .A0(n9750), .A1(n1256), .B0(n51), .B1(n1255), .C0(n1254), 
        .Y(stg2_real_Wn[51]) );
  OA22XL U975 ( .A0(n19), .A1(n2423), .B0(n197), .B1(n2965), .Y(n2422) );
  OA22XL U976 ( .A0(n9200), .A1(n2965), .B0(n19), .B1(n2508), .Y(n2507) );
  OA22XL U977 ( .A0(n45), .A1(n2428), .B0(n207), .B1(n2978), .Y(n2427) );
  OA22XL U978 ( .A0(n917), .A1(n2978), .B0(n48), .B1(n2514), .Y(n2513) );
  OA22XL U979 ( .A0(n906), .A1(n2978), .B0(n48), .B1(n2979), .Y(n2976) );
  OA22XL U980 ( .A0(n47), .A1(n2433), .B0(n183), .B1(n2991), .Y(n2432) );
  OA22XL U981 ( .A0(n9200), .A1(n2991), .B0(n45), .B1(n2520), .Y(n2519) );
  OA22XL U982 ( .A0(n20), .A1(n2438), .B0(n199), .B1(n3004), .Y(n2437) );
  OA22XL U983 ( .A0(n917), .A1(n3004), .B0(n46), .B1(n2526), .Y(n2525) );
  OA22XL U984 ( .A0(n917), .A1(n3017), .B0(n47), .B1(n2532), .Y(n2531) );
  OA22XL U985 ( .A0(n917), .A1(n3030), .B0(n49), .B1(n2538), .Y(n2537) );
  OA22XL U986 ( .A0(n917), .A1(n3043), .B0(n20), .B1(n2544), .Y(n2543) );
  OA22XL U987 ( .A0(n52), .A1(n2443), .B0(n187), .B1(n3017), .Y(n2442) );
  OA22XL U988 ( .A0(n46), .A1(n2448), .B0(n189), .B1(n3030), .Y(n2447) );
  OA22XL U989 ( .A0(n19), .A1(n2453), .B0(n195), .B1(n3043), .Y(n2452) );
  AOI2BB1XL U990 ( .A0N(n851), .A1N(n2636), .B0(n827), .Y(n2633) );
  AOI2BB1XL U991 ( .A0N(n851), .A1N(n2645), .B0(n828), .Y(n2642) );
  AOI2BB2XL U992 ( .B0(stg2_img_15__5_), .B1(n874), .A0N(n2991), .A1N(n852), 
        .Y(n2518) );
  AOI2BB1XL U993 ( .A0N(n851), .A1N(n2654), .B0(n829), .Y(n2651) );
  AOI2BB2XL U994 ( .B0(stg2_img_15__4_), .B1(n873), .A0N(n3004), .A1N(n852), 
        .Y(n2524) );
  OAI221XL U995 ( .A0(n9760), .A1(n2792), .B0(n50), .B1(n126), .C0(n1368), .Y(
        stg2_real_Wn[22]) );
  OAI221XL U996 ( .A0(n9760), .A1(n2782), .B0(n48), .B1(n125), .C0(n1360), .Y(
        stg2_real_Wn[23]) );
  OAI221XL U997 ( .A0(n9760), .A1(n2802), .B0(n52), .B1(n117), .C0(n1376), .Y(
        stg2_real_Wn[21]) );
  OAI221XL U998 ( .A0(n9770), .A1(n2804), .B0(n46), .B1(n2803), .C0(n2351), 
        .Y(stg2_real_Wn[37]) );
  OA22XL U999 ( .A0(n200), .A1(n2806), .B0(n78), .B1(n2350), .Y(n2351) );
  OAI221XL U1000 ( .A0(n9770), .A1(n2784), .B0(n52), .B1(n2783), .C0(n2337), 
        .Y(stg2_real_Wn[39]) );
  OA22XL U1001 ( .A0(n207), .A1(n2786), .B0(n84), .B1(n2336), .Y(n2337) );
  OAI221XL U1002 ( .A0(n9770), .A1(n2794), .B0(n20), .B1(n2793), .C0(n2344), 
        .Y(stg2_real_Wn[38]) );
  OA22XL U1003 ( .A0(n193), .A1(n2796), .B0(n79), .B1(n2343), .Y(n2344) );
  OAI221XL U1004 ( .A0(n9770), .A1(n2774), .B0(n50), .B1(n2773), .C0(n2330), 
        .Y(stg2_real_Wn[40]) );
  OA22XL U1005 ( .A0(n207), .A1(n2776), .B0(n75), .B1(n2329), .Y(n2330) );
  OAI221XL U1006 ( .A0(n9740), .A1(n2805), .B0(n50), .B1(n2801), .C0(n2650), 
        .Y(stg2_real_Wn[5]) );
  OAI221XL U1007 ( .A0(n9810), .A1(n2795), .B0(n48), .B1(n2791), .C0(n2641), 
        .Y(stg2_real_Wn[6]) );
  OAI221XL U1008 ( .A0(n9810), .A1(n2785), .B0(n46), .B1(n2781), .C0(n2632), 
        .Y(stg2_real_Wn[7]) );
  OAI221XL U1009 ( .A0(n9750), .A1(n1247), .B0(n48), .B1(n1246), .C0(n1245), 
        .Y(stg2_real_Wn[52]) );
  OAI221XL U1010 ( .A0(n9750), .A1(n1238), .B0(n45), .B1(n1237), .C0(n1236), 
        .Y(stg2_real_Wn[53]) );
  OAI221XL U1011 ( .A0(n9750), .A1(n1229), .B0(n19), .B1(n1228), .C0(n1227), 
        .Y(stg2_real_Wn[54]) );
  OAI221XL U1012 ( .A0(n9760), .A1(n2772), .B0(n46), .B1(n124), .C0(n1352), 
        .Y(stg2_real_Wn[24]) );
  OAI221XL U1013 ( .A0(n9760), .A1(n2762), .B0(n20), .B1(n1344), .C0(n1343), 
        .Y(stg2_real_Wn[25]) );
  OAI221XL U1014 ( .A0(n9760), .A1(n2752), .B0(n52), .B1(n1335), .C0(n1334), 
        .Y(stg2_real_Wn[26]) );
  OAI221XL U1015 ( .A0(n9770), .A1(n2764), .B0(n48), .B1(n2763), .C0(n2323), 
        .Y(stg2_real_Wn[41]) );
  OAI221XL U1016 ( .A0(n9770), .A1(n2754), .B0(n46), .B1(n2753), .C0(n2316), 
        .Y(stg2_real_Wn[42]) );
  OAI221XL U1017 ( .A0(n9770), .A1(n2744), .B0(n20), .B1(n2743), .C0(n2309), 
        .Y(stg2_real_Wn[43]) );
  OAI221XL U1018 ( .A0(n9800), .A1(n2775), .B0(n20), .B1(n2771), .C0(n2623), 
        .Y(stg2_real_Wn[8]) );
  OAI221XL U1019 ( .A0(n9800), .A1(n2765), .B0(n52), .B1(n2761), .C0(n2614), 
        .Y(stg2_real_Wn[9]) );
  OAI221XL U1020 ( .A0(n9800), .A1(n2755), .B0(n50), .B1(n2751), .C0(n2605), 
        .Y(stg2_real_Wn[10]) );
  OAI221XL U1021 ( .A0(n9740), .A1(n1220), .B0(n51), .B1(n1219), .C0(n1218), 
        .Y(stg2_real_Wn[55]) );
  OAI221XL U1022 ( .A0(n9740), .A1(n1211), .B0(n49), .B1(n1210), .C0(n1209), 
        .Y(stg2_real_Wn[56]) );
  OAI221XL U1023 ( .A0(n9740), .A1(n1202), .B0(n47), .B1(n1201), .C0(n1200), 
        .Y(stg2_real_Wn[57]) );
  OAI221XL U1024 ( .A0(n9740), .A1(n1193), .B0(n45), .B1(n1192), .C0(n1191), 
        .Y(stg2_real_Wn[58]) );
  OAI221XL U1025 ( .A0(n9750), .A1(n2732), .B0(n49), .B1(n1317), .C0(n1316), 
        .Y(stg2_real_Wn[28]) );
  OAI221XL U1026 ( .A0(n9750), .A1(n2722), .B0(n47), .B1(n1308), .C0(n1307), 
        .Y(stg2_real_Wn[29]) );
  OAI221XL U1027 ( .A0(n9750), .A1(n2742), .B0(n50), .B1(n1326), .C0(n1325), 
        .Y(stg2_real_Wn[27]) );
  OAI221XL U1028 ( .A0(n9770), .A1(n2724), .B0(n50), .B1(n2723), .C0(n1797), 
        .Y(stg2_real_Wn[45]) );
  OAI221XL U1029 ( .A0(n9770), .A1(n2714), .B0(n49), .B1(n92), .C0(n1434), .Y(
        stg2_real_Wn[46]) );
  OAI221XL U1030 ( .A0(n9770), .A1(n2734), .B0(n52), .B1(n2733), .C0(n1804), 
        .Y(stg2_real_Wn[44]) );
  OAI221XL U1031 ( .A0(n9740), .A1(n2745), .B0(n48), .B1(n2741), .C0(n2596), 
        .Y(stg2_real_Wn[11]) );
  OAI221XL U1032 ( .A0(n9790), .A1(n2735), .B0(n45), .B1(n2731), .C0(n2587), 
        .Y(stg2_real_Wn[12]) );
  OAI221XL U1033 ( .A0(n9740), .A1(n2725), .B0(n19), .B1(n2721), .C0(n2578), 
        .Y(stg2_real_Wn[13]) );
  OAI221XL U1034 ( .A0(n9790), .A1(n2715), .B0(n52), .B1(n2712), .C0(n2569), 
        .Y(stg2_real_Wn[14]) );
  OAI221XL U1035 ( .A0(n9740), .A1(n1184), .B0(n19), .B1(n1183), .C0(n1182), 
        .Y(stg2_real_Wn[59]) );
  OAI221XL U1036 ( .A0(n9740), .A1(n1175), .B0(n51), .B1(n1174), .C0(n1173), 
        .Y(stg2_real_Wn[60]) );
  OAI221XL U1037 ( .A0(n9740), .A1(n1166), .B0(n48), .B1(n1165), .C0(n1164), 
        .Y(stg2_real_Wn[61]) );
  INVXL U1038 ( .A(mul_2_Wn_19), .Y(n10520) );
  OAI221XL U1039 ( .A0(n9790), .A1(n3073), .B0(n47), .B1(n90), .C0(n2561), .Y(
        stg2_real_Wn[15]) );
  OAI221XL U1040 ( .A0(n9750), .A1(n89), .B0(n19), .B1(n152), .C0(n1291), .Y(
        stg2_real_Wn[31]) );
  OAI221XL U1041 ( .A0(n9750), .A1(n2713), .B0(n20), .B1(n1297), .C0(n1296), 
        .Y(stg2_real_Wn[30]) );
  OAI221XL U1042 ( .A0(n9740), .A1(n1157), .B0(n46), .B1(n1156), .C0(n1155), 
        .Y(stg2_real_Wn[62]) );
  OAI221XL U1043 ( .A0(n9800), .A1(n2707), .B0(n20), .B1(n2706), .C0(n2705), 
        .Y(stg2_real_Wn[63]) );
  OAI221XL U1044 ( .A0(n9760), .A1(n91), .B0(n50), .B1(n96), .C0(n1427), .Y(
        stg2_real_Wn[47]) );
  NAND3BXL U1045 ( .AN(n914), .B(n852), .C(n1300), .Y(n1284) );
  NAND2XL U1046 ( .A(n10480), .B(n10360), .Y(n7280) );
  NAND2XL U1047 ( .A(n791), .B(n10360), .Y(n7290) );
  OA22XL U1048 ( .A0(n78), .A1(n2984), .B0(n10350), .B1(n2983), .Y(n2985) );
  OA22XL U1049 ( .A0(n3120), .A1(n9280), .B0(n3072), .B1(n2980), .Y(n2987) );
  NAND4X4 U1050 ( .A(n179), .B(n2961), .C(n2960), .D(n2959), .Y(mul_1_in[8])
         );
  OA22XL U1051 ( .A0(n3111), .A1(n9280), .B0(n3072), .B1(n2954), .Y(n2961) );
  NAND4X4 U1052 ( .A(n2780), .B(n2779), .C(n2778), .D(n2777), .Y(mul_2_in[8])
         );
  OA22XL U1053 ( .A0(n49), .A1(n2774), .B0(n199), .B1(n2773), .Y(n2778) );
  OA22XL U1054 ( .A0(n3133), .A1(n9280), .B0(n9220), .B1(n3019), .Y(n3026) );
  OA22XL U1055 ( .A0(n3125), .A1(n9280), .B0(n3072), .B1(n2993), .Y(n3000) );
  OA22XL U1056 ( .A0(n82), .A1(n2997), .B0(n10460), .B1(n2996), .Y(n2998) );
  OA22XL U1057 ( .A0(n3141), .A1(n9280), .B0(n3072), .B1(n3045), .Y(n3052) );
  OA22XL U1058 ( .A0(n20), .A1(n2844), .B0(n9590), .B1(n2843), .Y(n2848) );
  OA22XL U1059 ( .A0(n76), .A1(n2846), .B0(n10350), .B1(n2845), .Y(n2847) );
  OA22XL U1060 ( .A0(n20), .A1(n3061), .B0(n187), .B1(n3060), .Y(n3065) );
  OA22XL U1061 ( .A0(n75), .A1(n3063), .B0(n10460), .B1(n3062), .Y(n3064) );
  OA22XL U1062 ( .A0(n49), .A1(n2917), .B0(n191), .B1(n2916), .Y(n2921) );
  OA22XL U1063 ( .A0(n80), .A1(n2919), .B0(n10460), .B1(n2918), .Y(n2920) );
  OA22XL U1064 ( .A0(n50), .A1(n2854), .B0(n9630), .B1(n2853), .Y(n2858) );
  OA22XL U1065 ( .A0(n84), .A1(n2856), .B0(n10350), .B1(n2855), .Y(n2857) );
  OA22XL U1066 ( .A0(n46), .A1(n2824), .B0(n205), .B1(n2823), .Y(n2828) );
  OA22XL U1067 ( .A0(n79), .A1(n2826), .B0(n10350), .B1(n2825), .Y(n2827) );
  OA22XL U1068 ( .A0(n45), .A1(n2804), .B0(n208), .B1(n2803), .Y(n2808) );
  OA22XL U1069 ( .A0(n79), .A1(n2806), .B0(n10350), .B1(n2805), .Y(n2807) );
  OA22XL U1070 ( .A0(n51), .A1(n2784), .B0(n181), .B1(n2783), .Y(n2788) );
  OA22XL U1071 ( .A0(n83), .A1(n2786), .B0(n10460), .B1(n2785), .Y(n2787) );
  INVX3 U1072 ( .A(n10450), .Y(n10530) );
  AND4XL U1073 ( .A(n1810), .B(n1811), .C(n177), .D(n176), .Y(n840) );
  AND2XL U1074 ( .A(n1790), .B(n1789), .Y(n838) );
  AOI222XL U1075 ( .A0(stg_reg[63]), .A1(n862), .B0(stg_reg[95]), .B1(n913), 
        .C0(n1728), .C1(n904), .Y(n3078) );
  AOI222XL U1076 ( .A0(stg_reg[47]), .A1(n861), .B0(n914), .B1(stg_reg[79]), 
        .C0(n904), .C1(n1552), .Y(n2874) );
  OA22XL U1077 ( .A0(n45), .A1(n2891), .B0(n195), .B1(n93), .Y(n2895) );
  OA22XL U1078 ( .A0(n75), .A1(n2893), .B0(n10460), .B1(n2892), .Y(n2894) );
  OA22XL U1079 ( .A0(n20), .A1(n110), .B0(n189), .B1(n95), .Y(n2883) );
  OA22XL U1080 ( .A0(n75), .A1(n2881), .B0(n10460), .B1(n2880), .Y(n2882) );
  OA22XL U1081 ( .A0(n51), .A1(n2714), .B0(n193), .B1(n92), .Y(n2718) );
  OA22XL U1082 ( .A0(n82), .A1(n2716), .B0(n10460), .B1(n2715), .Y(n2717) );
  OAI221XL U1083 ( .A0(n9740), .A1(n11410), .B0(n50), .B1(n11400), .C0(n11390), 
        .Y(stg2_img_Wn[49]) );
  OAI221XL U1084 ( .A0(n9740), .A1(n11350), .B0(n49), .B1(n11340), .C0(n11330), 
        .Y(stg2_img_Wn[50]) );
  OAI221XL U1085 ( .A0(n9740), .A1(n11290), .B0(n47), .B1(n11280), .C0(n11270), 
        .Y(stg2_img_Wn[51]) );
  OAI221XL U1086 ( .A0(n9780), .A1(n3047), .B0(n20), .B1(n3046), .C0(n2455), 
        .Y(stg2_img_Wn[33]) );
  OAI221XL U1087 ( .A0(n9780), .A1(n3034), .B0(n47), .B1(n3033), .C0(n2450), 
        .Y(stg2_img_Wn[34]) );
  OAI221XL U1088 ( .A0(n9780), .A1(n3021), .B0(n45), .B1(n3020), .C0(n2445), 
        .Y(stg2_img_Wn[35]) );
  OAI221XL U1089 ( .A0(n9760), .A1(n3137), .B0(n20), .B1(n99), .C0(n3136), .Y(
        stg2_img_Wn[18]) );
  OA22XL U1090 ( .A0(n9590), .A1(n3135), .B0(n76), .B1(n3134), .Y(n3136) );
  OAI221XL U1091 ( .A0(n9760), .A1(n3133), .B0(n19), .B1(n102), .C0(n3132), 
        .Y(stg2_img_Wn[19]) );
  OA22XL U1092 ( .A0(n193), .A1(n3131), .B0(n82), .B1(n3130), .Y(n3132) );
  OAI221XL U1093 ( .A0(n9790), .A1(n3048), .B0(n48), .B1(n3045), .C0(n2547), 
        .Y(stg2_img_Wn[1]) );
  OAI221XL U1094 ( .A0(n9790), .A1(n3035), .B0(n19), .B1(n3032), .C0(n2541), 
        .Y(stg2_img_Wn[2]) );
  OAI221XL U1095 ( .A0(n9790), .A1(n3022), .B0(n51), .B1(n3019), .C0(n2535), 
        .Y(stg2_img_Wn[3]) );
  OAI221XL U1096 ( .A0(n9760), .A1(n3141), .B0(n50), .B1(n100), .C0(n3140), 
        .Y(stg2_img_Wn[17]) );
  INVX1 U1097 ( .A(stg_reg[0]), .Y(n3062) );
  INVX1 U1098 ( .A(stg_reg[29]), .Y(n2725) );
  INVX1 U1099 ( .A(stg_reg[118]), .Y(n2796) );
  INVX1 U1100 ( .A(stg_reg[123]), .Y(n2746) );
  AO22XL U1101 ( .A0(stg_reg[142]), .A1(n843), .B0(stg4_img[62]), .B1(n209), 
        .Y(n2101) );
  AO22XL U1102 ( .A0(stg_reg[141]), .A1(n843), .B0(stg4_img[61]), .B1(n209), 
        .Y(n2102) );
  AO22XL U1103 ( .A0(stg_reg[143]), .A1(n843), .B0(stg4_img[63]), .B1(n209), 
        .Y(n2100) );
  OAI221XL U1104 ( .A0(n9750), .A1(n11230), .B0(n45), .B1(n11220), .C0(n11210), 
        .Y(stg2_img_Wn[52]) );
  OAI221XL U1105 ( .A0(n9750), .A1(n11170), .B0(n19), .B1(n11160), .C0(n11150), 
        .Y(stg2_img_Wn[53]) );
  OAI221XL U1106 ( .A0(n9810), .A1(n11110), .B0(n51), .B1(n11100), .C0(n11090), 
        .Y(stg2_img_Wn[54]) );
  OAI221XL U1107 ( .A0(n9780), .A1(n3008), .B0(n19), .B1(n3007), .C0(n2440), 
        .Y(stg2_img_Wn[36]) );
  OA22XL U1108 ( .A0(n189), .A1(n3010), .B0(n76), .B1(n2439), .Y(n2440) );
  OAI221XL U1109 ( .A0(n9780), .A1(n2995), .B0(n51), .B1(n2994), .C0(n2435), 
        .Y(stg2_img_Wn[37]) );
  OA22XL U1110 ( .A0(n187), .A1(n2997), .B0(n82), .B1(n2434), .Y(n2435) );
  OAI221XL U1111 ( .A0(n9780), .A1(n2982), .B0(n49), .B1(n2981), .C0(n2430), 
        .Y(stg2_img_Wn[38]) );
  OA22XL U1112 ( .A0(n202), .A1(n2984), .B0(n82), .B1(n2429), .Y(n2430) );
  OAI221XL U1113 ( .A0(n9760), .A1(n3129), .B0(n50), .B1(n101), .C0(n3128), 
        .Y(stg2_img_Wn[20]) );
  OA22XL U1114 ( .A0(n185), .A1(n3127), .B0(n84), .B1(n3126), .Y(n3128) );
  OAI221XL U1115 ( .A0(n9760), .A1(n3125), .B0(n49), .B1(n3124), .C0(n3123), 
        .Y(stg2_img_Wn[21]) );
  OA22XL U1116 ( .A0(n183), .A1(n3122), .B0(n81), .B1(n3121), .Y(n3123) );
  OAI221XL U1117 ( .A0(n9760), .A1(n3120), .B0(n47), .B1(n3119), .C0(n3118), 
        .Y(stg2_img_Wn[22]) );
  OA22XL U1118 ( .A0(n9590), .A1(n3117), .B0(n78), .B1(n3116), .Y(n3118) );
  OAI221XL U1119 ( .A0(n9790), .A1(n3009), .B0(n49), .B1(n3006), .C0(n2529), 
        .Y(stg2_img_Wn[4]) );
  OAI221XL U1120 ( .A0(n9790), .A1(n2996), .B0(n47), .B1(n2993), .C0(n2523), 
        .Y(stg2_img_Wn[5]) );
  OAI221XL U1121 ( .A0(n9790), .A1(n2983), .B0(n46), .B1(n2980), .C0(n2517), 
        .Y(stg2_img_Wn[6]) );
  AO22XL U1122 ( .A0(n1446), .A1(n9420), .B0(stg4_img[60]), .B1(n66), .Y(n2199) );
  AO22XL U1123 ( .A0(n1443), .A1(n9420), .B0(stg4_img[59]), .B1(n54), .Y(n2200) );
  AO22XL U1124 ( .A0(stg_reg[140]), .A1(n843), .B0(stg4_img[60]), .B1(n209), 
        .Y(n2103) );
  AO22XL U1125 ( .A0(stg_reg[139]), .A1(n843), .B0(stg4_img[59]), .B1(n209), 
        .Y(n2104) );
  AO22XL U1126 ( .A0(stg_reg[138]), .A1(n843), .B0(stg4_img[58]), .B1(n209), 
        .Y(n2105) );
  OAI221XL U1127 ( .A0(n9810), .A1(n11050), .B0(n49), .B1(n11040), .C0(n11030), 
        .Y(stg2_img_Wn[55]) );
  OAI221XL U1128 ( .A0(n9810), .A1(n10990), .B0(n47), .B1(n10980), .C0(n10970), 
        .Y(stg2_img_Wn[56]) );
  OAI221XL U1129 ( .A0(n9810), .A1(n10930), .B0(n45), .B1(n10920), .C0(n10910), 
        .Y(stg2_img_Wn[57]) );
  OAI221XL U1130 ( .A0(n9750), .A1(n2969), .B0(n47), .B1(n2968), .C0(n2425), 
        .Y(stg2_img_Wn[39]) );
  OA22XL U1131 ( .A0(n181), .A1(n2971), .B0(n77), .B1(n2424), .Y(n2425) );
  OAI221XL U1132 ( .A0(n9740), .A1(n2956), .B0(n45), .B1(n2955), .C0(n2420), 
        .Y(stg2_img_Wn[40]) );
  OA22XL U1133 ( .A0(n189), .A1(n2958), .B0(n78), .B1(n2419), .Y(n2420) );
  OAI221XL U1134 ( .A0(n9750), .A1(n2943), .B0(n19), .B1(n2942), .C0(n2415), 
        .Y(stg2_img_Wn[41]) );
  OA22XL U1135 ( .A0(n203), .A1(n2945), .B0(n84), .B1(n141), .Y(n2415) );
  OAI221XL U1136 ( .A0(n9750), .A1(n3115), .B0(n45), .B1(n105), .C0(n3114), 
        .Y(stg2_img_Wn[23]) );
  OAI221XL U1137 ( .A0(n9800), .A1(n3111), .B0(n19), .B1(n3110), .C0(n3109), 
        .Y(stg2_img_Wn[24]) );
  OA22XL U1138 ( .A0(n205), .A1(n3108), .B0(n84), .B1(n3107), .Y(n3109) );
  OAI221XL U1139 ( .A0(n9800), .A1(n3106), .B0(n51), .B1(n3105), .C0(n3104), 
        .Y(stg2_img_Wn[25]) );
  OAI221XL U1140 ( .A0(n9790), .A1(n2970), .B0(n20), .B1(n2967), .C0(n2511), 
        .Y(stg2_img_Wn[7]) );
  OAI221XL U1141 ( .A0(n9790), .A1(n2957), .B0(n52), .B1(n2954), .C0(n2505), 
        .Y(stg2_img_Wn[8]) );
  OAI221XL U1142 ( .A0(n9790), .A1(n2944), .B0(n50), .B1(n2941), .C0(n2499), 
        .Y(stg2_img_Wn[9]) );
  INVXL U1143 ( .A(stg_reg[64]), .Y(n3145) );
  INVXL U1144 ( .A(stg_reg[65]), .Y(n3139) );
  INVXL U1145 ( .A(stg_reg[32]), .Y(n2552) );
  INVXL U1146 ( .A(stg_reg[33]), .Y(n2546) );
  INVXL U1147 ( .A(stg_reg[80]), .Y(n1415) );
  INVXL U1148 ( .A(stg_reg[81]), .Y(n1407) );
  INVXL U1149 ( .A(stg_reg[82]), .Y(n1399) );
  INVXL U1150 ( .A(stg_reg[48]), .Y(n2696) );
  INVXL U1151 ( .A(stg_reg[49]), .Y(n2685) );
  INVXL U1152 ( .A(stg_reg[50]), .Y(n2676) );
  AO22XL U1153 ( .A0(stg_reg[137]), .A1(n843), .B0(stg4_img[57]), .B1(n209), 
        .Y(n2106) );
  AO22XL U1154 ( .A0(stg_reg[136]), .A1(n843), .B0(stg4_img[56]), .B1(n209), 
        .Y(n2107) );
  AO22XL U1155 ( .A0(stg_reg[135]), .A1(n843), .B0(stg4_img[55]), .B1(n209), 
        .Y(n2108) );
  OAI221XL U1156 ( .A0(n9760), .A1(n10880), .B0(n19), .B1(n10870), .C0(n10860), 
        .Y(stg2_img_Wn[58]) );
  OAI221XL U1157 ( .A0(n9800), .A1(n10830), .B0(n51), .B1(n10820), .C0(n10810), 
        .Y(stg2_img_Wn[59]) );
  OAI221XL U1158 ( .A0(n9810), .A1(n10780), .B0(n48), .B1(n10770), .C0(n10760), 
        .Y(stg2_img_Wn[60]) );
  OAI221XL U1159 ( .A0(n9740), .A1(n2930), .B0(n51), .B1(n2929), .C0(n2411), 
        .Y(stg2_img_Wn[42]) );
  OA22XL U1160 ( .A0(n193), .A1(n2932), .B0(n81), .B1(n142), .Y(n2411) );
  OAI221XL U1161 ( .A0(n9740), .A1(n2917), .B0(n49), .B1(n2916), .C0(n2407), 
        .Y(stg2_img_Wn[43]) );
  OA22XL U1162 ( .A0(n181), .A1(n2919), .B0(n83), .B1(n143), .Y(n2407) );
  OAI221XL U1163 ( .A0(n9820), .A1(n2904), .B0(n47), .B1(n2903), .C0(n2403), 
        .Y(stg2_img_Wn[44]) );
  OA22XL U1164 ( .A0(n205), .A1(n2906), .B0(n81), .B1(n144), .Y(n2403) );
  OAI221XL U1165 ( .A0(n9810), .A1(n2891), .B0(n45), .B1(n93), .C0(n2399), .Y(
        stg2_img_Wn[45]) );
  OAI221XL U1166 ( .A0(n9800), .A1(n3102), .B0(n49), .B1(n3101), .C0(n3100), 
        .Y(stg2_img_Wn[26]) );
  OAI221XL U1167 ( .A0(n9800), .A1(n3098), .B0(n47), .B1(n3097), .C0(n3096), 
        .Y(stg2_img_Wn[27]) );
  OAI221XL U1168 ( .A0(n9790), .A1(n2931), .B0(n48), .B1(n2928), .C0(n2494), 
        .Y(stg2_img_Wn[10]) );
  OAI221XL U1169 ( .A0(n9780), .A1(n2918), .B0(n46), .B1(n2915), .C0(n2489), 
        .Y(stg2_img_Wn[11]) );
  OAI221XL U1170 ( .A0(n9780), .A1(n2905), .B0(n20), .B1(n2902), .C0(n2484), 
        .Y(stg2_img_Wn[12]) );
  OAI221XL U1171 ( .A0(n9780), .A1(n2892), .B0(n52), .B1(n108), .C0(n2479), 
        .Y(stg2_img_Wn[13]) );
  OAI221XL U1172 ( .A0(n9800), .A1(n3094), .B0(n46), .B1(n3093), .C0(n3092), 
        .Y(stg2_img_Wn[28]) );
  OAI221XL U1173 ( .A0(n9800), .A1(n3090), .B0(n20), .B1(n132), .C0(n3089), 
        .Y(stg2_img_Wn[29]) );
  INVXL U1174 ( .A(stg_reg[66]), .Y(n3135) );
  INVXL U1175 ( .A(stg_reg[67]), .Y(n3131) );
  INVXL U1176 ( .A(stg_reg[68]), .Y(n3127) );
  INVXL U1177 ( .A(stg_reg[34]), .Y(n2540) );
  INVXL U1178 ( .A(stg_reg[35]), .Y(n2534) );
  INVXL U1179 ( .A(stg_reg[36]), .Y(n2528) );
  INVXL U1180 ( .A(stg_reg[83]), .Y(n1391) );
  INVXL U1181 ( .A(stg_reg[84]), .Y(n1383) );
  INVXL U1182 ( .A(stg_reg[85]), .Y(n1375) );
  INVXL U1183 ( .A(stg_reg[51]), .Y(n2667) );
  INVXL U1184 ( .A(stg_reg[52]), .Y(n2658) );
  INVXL U1185 ( .A(stg_reg[53]), .Y(n2649) );
  AO22XL U1186 ( .A0(stg_reg[134]), .A1(n843), .B0(stg4_img[54]), .B1(n209), 
        .Y(n2109) );
  AO22XL U1187 ( .A0(stg_reg[133]), .A1(n843), .B0(stg4_img[53]), .B1(n209), 
        .Y(n2110) );
  AO22XL U1188 ( .A0(stg_reg[132]), .A1(n843), .B0(stg4_img[52]), .B1(n209), 
        .Y(n2111) );
  OAI221XL U1189 ( .A0(n9770), .A1(n10730), .B0(n46), .B1(n10720), .C0(n10710), 
        .Y(stg2_img_Wn[61]) );
  OAI221XL U1190 ( .A0(n9770), .A1(n10680), .B0(n45), .B1(n10670), .C0(n10660), 
        .Y(stg2_img_Wn[62]) );
  OAI221XL U1191 ( .A0(n9780), .A1(n2869), .B0(n52), .B1(n111), .C0(n2469), 
        .Y(stg2_img_Wn[15]) );
  OAI221XL U1192 ( .A0(n9800), .A1(n97), .B0(n48), .B1(n150), .C0(n3085), .Y(
        stg2_img_Wn[31]) );
  OAI221XL U1193 ( .A0(n9820), .A1(n110), .B0(n19), .B1(n95), .C0(n2395), .Y(
        stg2_img_Wn[46]) );
  OAI221XL U1194 ( .A0(n9780), .A1(n2880), .B0(n50), .B1(n112), .C0(n2474), 
        .Y(stg2_img_Wn[14]) );
  OAI221XL U1195 ( .A0(n9800), .A1(n94), .B0(n51), .B1(n151), .C0(n3087), .Y(
        stg2_img_Wn[30]) );
  OAI221XL U1196 ( .A0(n9750), .A1(n10630), .B0(n49), .B1(n10620), .C0(n10610), 
        .Y(stg2_img_Wn[63]) );
  OAI221XL U1197 ( .A0(n9810), .A1(n113), .B0(n51), .B1(n2868), .C0(n2391), 
        .Y(stg2_img_Wn[47]) );
  OA22XL U1198 ( .A0(n205), .A1(n2870), .B0(n81), .B1(n171), .Y(n2391) );
  INVXL U1199 ( .A(stg_reg[69]), .Y(n3122) );
  INVXL U1200 ( .A(stg_reg[70]), .Y(n3117) );
  INVXL U1201 ( .A(stg_reg[71]), .Y(n3113) );
  INVXL U1202 ( .A(stg_reg[72]), .Y(n3108) );
  INVXL U1203 ( .A(stg_reg[37]), .Y(n2522) );
  INVXL U1204 ( .A(stg_reg[38]), .Y(n2516) );
  INVXL U1205 ( .A(stg_reg[39]), .Y(n2510) );
  INVXL U1206 ( .A(stg_reg[40]), .Y(n2504) );
  INVXL U1207 ( .A(stg_reg[86]), .Y(n1367) );
  INVXL U1208 ( .A(stg_reg[87]), .Y(n1359) );
  INVXL U1209 ( .A(stg_reg[88]), .Y(n1351) );
  INVXL U1210 ( .A(stg_reg[54]), .Y(n2640) );
  INVXL U1211 ( .A(stg_reg[55]), .Y(n2631) );
  INVXL U1212 ( .A(stg_reg[56]), .Y(n2622) );
  INVXL U1213 ( .A(stg_reg[57]), .Y(n2613) );
  AO22XL U1214 ( .A0(stg_reg[131]), .A1(n843), .B0(stg4_img[51]), .B1(n209), 
        .Y(n2112) );
  AO22XL U1215 ( .A0(stg_reg[130]), .A1(n843), .B0(stg4_img[50]), .B1(n209), 
        .Y(n2113) );
  AO22XL U1216 ( .A0(stg_reg[129]), .A1(n843), .B0(stg4_img[49]), .B1(n209), 
        .Y(n2114) );
  NAND2XL U1217 ( .A(n10510), .B(n10500), .Y(n1300) );
  MX2XL U1218 ( .A(n10360), .B(n10490), .S0(n1811), .Y(n10510) );
  AND2XL U1219 ( .A(n176), .B(n10360), .Y(n10490) );
  INVXL U1220 ( .A(stg_reg[73]), .Y(n3103) );
  INVXL U1221 ( .A(stg_reg[74]), .Y(n3099) );
  INVXL U1222 ( .A(stg_reg[75]), .Y(n3095) );
  INVXL U1223 ( .A(stg_reg[41]), .Y(n2498) );
  INVXL U1224 ( .A(stg_reg[42]), .Y(n2493) );
  INVXL U1225 ( .A(stg_reg[43]), .Y(n2488) );
  INVXL U1226 ( .A(stg_reg[89]), .Y(n1342) );
  INVXL U1227 ( .A(stg_reg[90]), .Y(n1333) );
  INVXL U1228 ( .A(stg_reg[91]), .Y(n1324) );
  INVXL U1229 ( .A(stg_reg[58]), .Y(n2604) );
  AO22XL U1230 ( .A0(stg_reg[128]), .A1(n843), .B0(stg4_img[48]), .B1(n209), 
        .Y(n2115) );
  INVXL U1231 ( .A(stg_reg[76]), .Y(n3091) );
  INVXL U1232 ( .A(stg_reg[92]), .Y(n1315) );
  AOI2BB1XL U1233 ( .A0N(n1811), .A1N(n1789), .B0(n176), .Y(n10390) );
  NAND2XL U1234 ( .A(n10360), .B(n10500), .Y(n10410) );
  AND2XL U1235 ( .A(fir_valid), .B(n1789), .Y(n842) );
  MX2XL U1236 ( .A(n842), .B(n10380), .S0(n1811), .Y(N36) );
  INVX3 U1237 ( .A(n3142), .Y(n9380) );
  INVX3 U1238 ( .A(n9470), .Y(n9360) );
  INVX3 U1239 ( .A(n9470), .Y(n9370) );
  INVX3 U1240 ( .A(n9470), .Y(n9390) );
  INVX3 U1241 ( .A(n9470), .Y(n9400) );
  INVX3 U1242 ( .A(mul_o_add[26]), .Y(n2926) );
  INVX3 U1243 ( .A(mul_o_add[24]), .Y(n2952) );
  INVX3 U1244 ( .A(mul_o_sub[26]), .Y(n2600) );
  INVX3 U1245 ( .A(mul_o_sub[24]), .Y(n2618) );
  INVX3 U1246 ( .A(mul_o_sub[29]), .Y(n2573) );
  INVX3 U1247 ( .A(mul_o_sub[25]), .Y(n2609) );
  INVX3 U1248 ( .A(mul_o_sub[23]), .Y(n2627) );
  INVX3 U1249 ( .A(mul_o_add[29]), .Y(n2889) );
  INVX3 U1250 ( .A(mul_o_add[25]), .Y(n2939) );
  INVX3 U1251 ( .A(mul_o_add[22]), .Y(n2978) );
  INVX3 U1252 ( .A(mul_o_add[20]), .Y(n3004) );
  INVX3 U1253 ( .A(mul_o_add[18]), .Y(n3030) );
  INVX3 U1254 ( .A(mul_o_sub[22]), .Y(n2636) );
  INVX3 U1255 ( .A(mul_o_sub[20]), .Y(n2654) );
  INVX3 U1256 ( .A(mul_o_sub[18]), .Y(n2672) );
  INVX3 U1257 ( .A(mul_o_sub[21]), .Y(n2645) );
  INVX3 U1258 ( .A(mul_o_sub[17]), .Y(n2681) );
  INVX3 U1259 ( .A(mul_o_add[23]), .Y(n2965) );
  INVX3 U1260 ( .A(mul_o_add[21]), .Y(n2991) );
  INVX3 U1261 ( .A(mul_o_add[19]), .Y(n3017) );
  INVX3 U1262 ( .A(mul_o_add[17]), .Y(n3043) );
  INVX3 U1263 ( .A(mul_o_add[16]), .Y(n3057) );
  INVX3 U1264 ( .A(mul_o_sub[16]), .Y(n2692) );
  CLKBUFX3 U1265 ( .A(n9470), .Y(n9440) );
  CLKBUFX3 U1266 ( .A(n9470), .Y(n9450) );
  CLKBUFX3 U1267 ( .A(n9470), .Y(n9410) );
  CLKBUFX3 U1268 ( .A(n9470), .Y(n9460) );
  CLKBUFX3 U1269 ( .A(n9470), .Y(n9420) );
  CLKBUFX3 U1270 ( .A(n9470), .Y(n9430) );
  INVX3 U1271 ( .A(mul_o_add[28]), .Y(n2900) );
  INVX3 U1272 ( .A(mul_o_sub[28]), .Y(n2582) );
  INVX3 U1273 ( .A(mul_o_sub[27]), .Y(n2591) );
  INVX3 U1274 ( .A(mul_o_add[27]), .Y(n2913) );
  INVX3 U1275 ( .A(mul_o_add[31]), .Y(n3081) );
  CLKBUFX3 U1276 ( .A(n9810), .Y(n9740) );
  CLKBUFX3 U1277 ( .A(n9820), .Y(n9790) );
  CLKBUFX3 U1278 ( .A(n9810), .Y(n9750) );
  CLKBUFX3 U1279 ( .A(n3142), .Y(n9470) );
  INVX3 U1280 ( .A(n10170), .Y(n9890) );
  INVX3 U1281 ( .A(n10150), .Y(n9940) );
  INVX3 U1282 ( .A(n10140), .Y(n9990) );
  INVX3 U1283 ( .A(n10120), .Y(n10040) );
  INVX3 U1284 ( .A(n10180), .Y(n9870) );
  INVX3 U1285 ( .A(n10160), .Y(n9920) );
  INVX3 U1286 ( .A(n10140), .Y(n9970) );
  INVX3 U1287 ( .A(n10130), .Y(n10020) );
  INVX3 U1288 ( .A(n10110), .Y(n10070) );
  INVX3 U1289 ( .A(n10180), .Y(n9850) );
  INVX3 U1290 ( .A(n10170), .Y(n9900) );
  INVX3 U1291 ( .A(n10150), .Y(n9950) );
  INVX3 U1292 ( .A(n10130), .Y(n10000) );
  INVX3 U1293 ( .A(n10120), .Y(n10050) );
  INVX3 U1294 ( .A(n10110), .Y(n10080) );
  INVX3 U1295 ( .A(n10110), .Y(n10060) );
  INVX3 U1296 ( .A(n10120), .Y(n10030) );
  INVX3 U1297 ( .A(n10130), .Y(n10010) );
  INVX3 U1298 ( .A(n10140), .Y(n9980) );
  INVX3 U1299 ( .A(n10150), .Y(n9960) );
  INVX3 U1300 ( .A(n10160), .Y(n9930) );
  INVX3 U1301 ( .A(n10160), .Y(n9910) );
  INVX3 U1302 ( .A(n10170), .Y(n9880) );
  INVX3 U1303 ( .A(n10180), .Y(n9860) );
  INVX3 U1304 ( .A(n10190), .Y(n9840) );
  CLKINVX1 U1305 ( .A(mul_2_Wn_11), .Y(n10440) );
  CLKINVX1 U1306 ( .A(mul_0_Wn[15]), .Y(n10540) );
  CLKBUFX3 U1307 ( .A(n7310), .Y(n856) );
  CLKBUFX3 U1308 ( .A(n2700), .Y(n844) );
  CLKINVX1 U1309 ( .A(n843), .Y(n2700) );
  INVX3 U1310 ( .A(n868), .Y(n883) );
  INVX3 U1311 ( .A(n887), .Y(n879) );
  INVX3 U1312 ( .A(n868), .Y(n882) );
  INVX3 U1313 ( .A(n868), .Y(n881) );
  INVX3 U1314 ( .A(n887), .Y(n880) );
  INVX3 U1315 ( .A(n868), .Y(n884) );
  INVX3 U1316 ( .A(n868), .Y(n878) );
  INVX3 U1317 ( .A(n868), .Y(n885) );
  CLKBUFX3 U1318 ( .A(n7310), .Y(n855) );
  INVX3 U1319 ( .A(n868), .Y(n886) );
  CLKBUFX3 U1320 ( .A(n9830), .Y(n10180) );
  CLKBUFX3 U1321 ( .A(n9830), .Y(n10170) );
  CLKBUFX3 U1322 ( .A(n9830), .Y(n10160) );
  CLKBUFX3 U1323 ( .A(n9830), .Y(n10150) );
  CLKBUFX3 U1324 ( .A(n9830), .Y(n10140) );
  CLKBUFX3 U1325 ( .A(n9830), .Y(n10130) );
  CLKBUFX3 U1326 ( .A(n9830), .Y(n10120) );
  CLKBUFX3 U1327 ( .A(n9830), .Y(n10110) );
  CLKBUFX3 U1328 ( .A(n7290), .Y(n10190) );
  INVX3 U1329 ( .A(n899), .Y(n873) );
  INVX3 U1330 ( .A(n900), .Y(n874) );
  INVX3 U1331 ( .A(n887), .Y(n875) );
  INVX3 U1332 ( .A(n899), .Y(n869) );
  INVX3 U1333 ( .A(n899), .Y(n870) );
  INVX3 U1334 ( .A(n887), .Y(n872) );
  INVX3 U1335 ( .A(n900), .Y(n871) );
  INVX3 U1336 ( .A(n900), .Y(n877) );
  INVX3 U1337 ( .A(n887), .Y(n876) );
  CLKBUFX3 U1338 ( .A(n10340), .Y(n10310) );
  CLKBUFX3 U1339 ( .A(n10340), .Y(n10300) );
  CLKBUFX3 U1340 ( .A(n10340), .Y(n10290) );
  CLKBUFX3 U1341 ( .A(n10340), .Y(n10280) );
  CLKBUFX3 U1342 ( .A(n10340), .Y(n10270) );
  CLKBUFX3 U1343 ( .A(n10190), .Y(n10250) );
  CLKBUFX3 U1344 ( .A(n10190), .Y(n10240) );
  CLKBUFX3 U1345 ( .A(n10190), .Y(n10230) );
  CLKBUFX3 U1346 ( .A(n10190), .Y(n10220) );
  CLKBUFX3 U1347 ( .A(n10190), .Y(n10210) );
  CLKBUFX3 U1348 ( .A(n10340), .Y(n10200) );
  CLKBUFX3 U1349 ( .A(n10340), .Y(n10260) );
  INVX3 U1350 ( .A(n9830), .Y(n10090) );
  INVX3 U1351 ( .A(n9830), .Y(n10100) );
  NAND2X1 U1352 ( .A(n7320), .B(n2865), .Y(mul_0_Wn_8) );
  INVX3 U1353 ( .A(n863), .Y(n861) );
  INVX3 U1354 ( .A(n863), .Y(n862) );
  CLKINVX1 U1355 ( .A(stg4_real[62]), .Y(n1152) );
  CLKINVX1 U1356 ( .A(stg4_real[61]), .Y(n1161) );
  CLKINVX1 U1357 ( .A(stg4_real[60]), .Y(n1170) );
  CLKINVX1 U1358 ( .A(stg4_real[59]), .Y(n1179) );
  CLKINVX1 U1359 ( .A(stg4_real[58]), .Y(n1188) );
  CLKINVX1 U1360 ( .A(stg4_real[57]), .Y(n1197) );
  CLKINVX1 U1361 ( .A(stg4_real[56]), .Y(n1206) );
  CLKINVX1 U1362 ( .A(stg4_real[46]), .Y(n1432) );
  CLKINVX1 U1363 ( .A(stg4_real[45]), .Y(n1795) );
  CLKINVX1 U1364 ( .A(stg4_real[44]), .Y(n1802) );
  CLKINVX1 U1365 ( .A(stg4_real[43]), .Y(n1809) );
  CLKINVX1 U1366 ( .A(stg4_real[42]), .Y(n2314) );
  CLKINVX1 U1367 ( .A(stg4_real[41]), .Y(n2321) );
  CLKINVX1 U1368 ( .A(stg4_real[40]), .Y(n2328) );
  CLKINVX1 U1369 ( .A(stg4_real[55]), .Y(n1215) );
  CLKINVX1 U1370 ( .A(stg4_real[54]), .Y(n1224) );
  CLKINVX1 U1371 ( .A(stg4_real[53]), .Y(n1233) );
  CLKINVX1 U1372 ( .A(stg4_real[52]), .Y(n1242) );
  CLKINVX1 U1373 ( .A(stg4_real[51]), .Y(n1251) );
  CLKINVX1 U1374 ( .A(stg4_real[50]), .Y(n1260) );
  CLKINVX1 U1375 ( .A(stg4_real[49]), .Y(n1269) );
  CLKINVX1 U1376 ( .A(stg4_real[39]), .Y(n2335) );
  CLKINVX1 U1377 ( .A(stg4_real[38]), .Y(n2342) );
  CLKINVX1 U1378 ( .A(stg4_real[37]), .Y(n2349) );
  CLKINVX1 U1379 ( .A(stg4_real[36]), .Y(n2356) );
  CLKINVX1 U1380 ( .A(stg4_real[35]), .Y(n2363) );
  CLKINVX1 U1381 ( .A(stg4_real[34]), .Y(n2370) );
  CLKINVX1 U1382 ( .A(stg4_real[33]), .Y(n2377) );
  CLKBUFX3 U1383 ( .A(n7330), .Y(n860) );
  CLKBUFX3 U1384 ( .A(n7340), .Y(n859) );
  CLKBUFX3 U1385 ( .A(n3079), .Y(n9240) );
  CLKBUFX3 U1386 ( .A(n3079), .Y(n9230) );
  CLKINVX1 U1387 ( .A(n10570), .Y(n1301) );
  NAND3BX1 U1388 ( .AN(n10560), .B(n7320), .C(n9340), .Y(n10570) );
  CLKBUFX3 U1389 ( .A(n1149), .Y(n843) );
  NAND2X1 U1390 ( .A(n858), .B(n866), .Y(n1149) );
  CLKBUFX3 U1391 ( .A(n2460), .Y(n850) );
  CLKBUFX3 U1392 ( .A(n2458), .Y(n848) );
  CLKBUFX3 U1393 ( .A(n107), .Y(n902) );
  CLKBUFX3 U1394 ( .A(n2458), .Y(n847) );
  CLKBUFX3 U1395 ( .A(n107), .Y(n901) );
  CLKBUFX3 U1396 ( .A(n2460), .Y(n849) );
  CLKBUFX3 U1397 ( .A(n9350), .Y(n9340) );
  CLKBUFX3 U1398 ( .A(n2456), .Y(n846) );
  CLKBUFX3 U1399 ( .A(n2456), .Y(n845) );
  CLKBUFX3 U1400 ( .A(n868), .Y(n887) );
  CLKBUFX3 U1401 ( .A(n893), .Y(n888) );
  CLKBUFX3 U1402 ( .A(n900), .Y(n892) );
  CLKBUFX3 U1403 ( .A(n900), .Y(n891) );
  CLKBUFX3 U1404 ( .A(n892), .Y(n889) );
  CLKBUFX3 U1405 ( .A(n894), .Y(n890) );
  CLKBUFX3 U1406 ( .A(n899), .Y(n895) );
  CLKBUFX3 U1407 ( .A(n900), .Y(n894) );
  CLKBUFX3 U1408 ( .A(n900), .Y(n893) );
  CLKBUFX3 U1409 ( .A(n9280), .Y(n9270) );
  CLKBUFX3 U1410 ( .A(n899), .Y(n896) );
  CLKBUFX3 U1411 ( .A(n899), .Y(n897) );
  CLKBUFX3 U1412 ( .A(n9280), .Y(n9260) );
  CLKBUFX3 U1413 ( .A(n899), .Y(n898) );
  CLKBUFX3 U1414 ( .A(n9330), .Y(n9310) );
  CLKBUFX3 U1415 ( .A(n9330), .Y(n9320) );
  CLKBUFX3 U1416 ( .A(n9350), .Y(n9330) );
  CLKBUFX3 U1417 ( .A(n9830), .Y(n10340) );
  NAND2X1 U1418 ( .A(n915), .B(n10470), .Y(mul_2_Wn_19) );
  CLKBUFX3 U1419 ( .A(n3082), .Y(n9250) );
  CLKINVX1 U1420 ( .A(stg4_img[15]), .Y(n2467) );
  CLKINVX1 U1421 ( .A(stg4_img[47]), .Y(n2390) );
  CLKINVX1 U1422 ( .A(stg4_real[63]), .Y(n2702) );
  CLKINVX1 U1423 ( .A(stg4_real[30]), .Y(n2710) );
  CLKINVX1 U1424 ( .A(stg4_real[29]), .Y(n1304) );
  CLKINVX1 U1425 ( .A(stg4_real[28]), .Y(n1313) );
  CLKINVX1 U1426 ( .A(stg4_real[27]), .Y(n1322) );
  CLKINVX1 U1427 ( .A(stg4_real[26]), .Y(n1331) );
  CLKINVX1 U1428 ( .A(stg4_real[25]), .Y(n1340) );
  CLKINVX1 U1429 ( .A(stg4_real[24]), .Y(n1349) );
  CLKINVX1 U1430 ( .A(stg4_real[14]), .Y(n2566) );
  CLKINVX1 U1431 ( .A(stg4_real[13]), .Y(n2575) );
  CLKINVX1 U1432 ( .A(stg4_real[12]), .Y(n2584) );
  CLKINVX1 U1433 ( .A(stg4_real[11]), .Y(n2593) );
  CLKINVX1 U1434 ( .A(stg4_real[10]), .Y(n2602) );
  CLKINVX1 U1435 ( .A(stg4_real[9]), .Y(n2611) );
  CLKINVX1 U1436 ( .A(stg4_real[8]), .Y(n2620) );
  CLKINVX1 U1437 ( .A(stg4_img[13]), .Y(n2477) );
  CLKINVX1 U1438 ( .A(stg4_img[12]), .Y(n2482) );
  CLKINVX1 U1439 ( .A(stg4_img[11]), .Y(n2487) );
  CLKINVX1 U1440 ( .A(stg4_img[10]), .Y(n2492) );
  CLKINVX1 U1441 ( .A(stg4_img[9]), .Y(n2497) );
  CLKINVX1 U1442 ( .A(stg4_img[8]), .Y(n2502) );
  CLKINVX1 U1443 ( .A(stg4_img[7]), .Y(n2508) );
  CLKINVX1 U1444 ( .A(stg4_img[29]), .Y(n2890) );
  CLKINVX1 U1445 ( .A(stg4_img[28]), .Y(n2901) );
  CLKINVX1 U1446 ( .A(stg4_img[27]), .Y(n2914) );
  CLKINVX1 U1447 ( .A(stg4_img[26]), .Y(n2927) );
  CLKINVX1 U1448 ( .A(stg4_img[25]), .Y(n2940) );
  CLKINVX1 U1449 ( .A(stg4_img[24]), .Y(n2953) );
  CLKINVX1 U1450 ( .A(stg4_img[46]), .Y(n2394) );
  CLKINVX1 U1451 ( .A(stg4_img[45]), .Y(n2398) );
  CLKINVX1 U1452 ( .A(stg4_img[44]), .Y(n2402) );
  CLKINVX1 U1453 ( .A(stg4_img[43]), .Y(n2406) );
  CLKINVX1 U1454 ( .A(stg4_img[42]), .Y(n2410) );
  CLKINVX1 U1455 ( .A(stg4_img[41]), .Y(n2414) );
  CLKINVX1 U1456 ( .A(stg4_img[40]), .Y(n2418) );
  CLKINVX1 U1457 ( .A(stg4_img[63]), .Y(n10550) );
  CLKINVX1 U1458 ( .A(stg4_img[62]), .Y(n10640) );
  CLKINVX1 U1459 ( .A(stg4_img[61]), .Y(n10690) );
  CLKINVX1 U1460 ( .A(stg4_img[60]), .Y(n10740) );
  CLKINVX1 U1461 ( .A(stg4_img[59]), .Y(n10790) );
  CLKINVX1 U1462 ( .A(stg4_img[58]), .Y(n10840) );
  CLKINVX1 U1463 ( .A(stg4_img[57]), .Y(n10890) );
  CLKINVX1 U1464 ( .A(stg4_real[47]), .Y(n1425) );
  AND2X2 U1465 ( .A(n856), .B(n9200), .Y(n7330) );
  AND2X2 U1466 ( .A(n854), .B(n852), .Y(n7340) );
  CLKINVX1 U1467 ( .A(stg4_real[23]), .Y(n1357) );
  CLKINVX1 U1468 ( .A(stg4_real[22]), .Y(n1365) );
  CLKINVX1 U1469 ( .A(stg4_real[21]), .Y(n1373) );
  CLKINVX1 U1470 ( .A(stg4_real[20]), .Y(n1381) );
  CLKINVX1 U1471 ( .A(stg4_real[19]), .Y(n1389) );
  CLKINVX1 U1472 ( .A(stg4_real[18]), .Y(n1397) );
  CLKINVX1 U1473 ( .A(stg4_real[17]), .Y(n1405) );
  CLKINVX1 U1474 ( .A(stg4_real[7]), .Y(n2629) );
  CLKINVX1 U1475 ( .A(stg4_real[6]), .Y(n2638) );
  CLKINVX1 U1476 ( .A(stg4_real[5]), .Y(n2647) );
  CLKINVX1 U1477 ( .A(stg4_real[4]), .Y(n2656) );
  CLKINVX1 U1478 ( .A(stg4_real[3]), .Y(n2665) );
  CLKINVX1 U1479 ( .A(stg4_real[2]), .Y(n2674) );
  CLKINVX1 U1480 ( .A(stg4_real[1]), .Y(n2683) );
  CLKINVX1 U1481 ( .A(stg4_real[0]), .Y(n2694) );
  CLKINVX1 U1482 ( .A(stg4_real[32]), .Y(n2384) );
  CLKINVX1 U1483 ( .A(stg4_real[48]), .Y(n1278) );
  CLKINVX1 U1484 ( .A(stg4_img[0]), .Y(n2550) );
  CLKINVX1 U1485 ( .A(stg4_img[16]), .Y(n3058) );
  CLKINVX1 U1486 ( .A(stg4_img[32]), .Y(n2461) );
  CLKINVX1 U1487 ( .A(stg4_img[6]), .Y(n2514) );
  CLKINVX1 U1488 ( .A(stg4_img[5]), .Y(n2520) );
  CLKINVX1 U1489 ( .A(stg4_img[4]), .Y(n2526) );
  CLKINVX1 U1490 ( .A(stg4_img[3]), .Y(n2532) );
  CLKINVX1 U1491 ( .A(stg4_img[2]), .Y(n2538) );
  CLKINVX1 U1492 ( .A(stg4_img[1]), .Y(n2544) );
  CLKINVX1 U1493 ( .A(stg4_img[23]), .Y(n2966) );
  CLKINVX1 U1494 ( .A(stg4_img[22]), .Y(n2979) );
  CLKINVX1 U1495 ( .A(stg4_img[21]), .Y(n2992) );
  CLKINVX1 U1496 ( .A(stg4_img[20]), .Y(n3005) );
  CLKINVX1 U1497 ( .A(stg4_img[19]), .Y(n3018) );
  CLKINVX1 U1498 ( .A(stg4_img[18]), .Y(n3031) );
  CLKINVX1 U1499 ( .A(stg4_img[17]), .Y(n3044) );
  CLKINVX1 U1500 ( .A(stg4_img[39]), .Y(n2423) );
  CLKINVX1 U1501 ( .A(stg4_img[38]), .Y(n2428) );
  CLKINVX1 U1502 ( .A(stg4_img[37]), .Y(n2433) );
  CLKINVX1 U1503 ( .A(stg4_img[36]), .Y(n2438) );
  CLKINVX1 U1504 ( .A(stg4_img[35]), .Y(n2443) );
  CLKINVX1 U1505 ( .A(stg4_img[34]), .Y(n2448) );
  CLKINVX1 U1506 ( .A(stg4_img[33]), .Y(n2453) );
  CLKINVX1 U1507 ( .A(stg4_img[48]), .Y(n11420) );
  CLKINVX1 U1508 ( .A(stg4_img[56]), .Y(n10940) );
  CLKINVX1 U1509 ( .A(stg4_img[55]), .Y(n11000) );
  CLKINVX1 U1510 ( .A(stg4_img[54]), .Y(n11060) );
  CLKINVX1 U1511 ( .A(stg4_img[53]), .Y(n11120) );
  CLKINVX1 U1512 ( .A(stg4_img[52]), .Y(n11180) );
  CLKINVX1 U1513 ( .A(stg4_img[51]), .Y(n11240) );
  CLKINVX1 U1514 ( .A(stg4_img[50]), .Y(n11300) );
  CLKINVX1 U1515 ( .A(stg4_img[49]), .Y(n11360) );
  CLKINVX1 U1516 ( .A(n1420), .Y(n1287) );
  CLKBUFX3 U1517 ( .A(n2690), .Y(n858) );
  CLKBUFX3 U1518 ( .A(n2690), .Y(n857) );
  CLKBUFX3 U1519 ( .A(n851), .Y(n852) );
  CLKBUFX3 U1520 ( .A(n9290), .Y(n9350) );
  CLKBUFX3 U1521 ( .A(n9330), .Y(n9300) );
  CLKBUFX3 U1522 ( .A(n10340), .Y(n10330) );
  CLKBUFX3 U1523 ( .A(n10340), .Y(n10320) );
  CLKBUFX3 U1524 ( .A(n868), .Y(n899) );
  CLKBUFX3 U1525 ( .A(n868), .Y(n900) );
  NAND2X1 U1526 ( .A(n2864), .B(n10460), .Y(mul_2_Wn_8) );
  CLKINVX1 U1527 ( .A(stg4_real[15]), .Y(n2558) );
  AND2X2 U1528 ( .A(n3205), .B(n7470), .Y(n7350) );
  AND2X2 U1529 ( .A(n3206), .B(n7350), .Y(n7360) );
  AND2X2 U1530 ( .A(n3207), .B(n7360), .Y(n7370) );
  AND2X2 U1531 ( .A(n3195), .B(n3194), .Y(n7380) );
  AND2X2 U1532 ( .A(n3196), .B(n7380), .Y(n7390) );
  AND2X2 U1533 ( .A(n3197), .B(n7390), .Y(n7400) );
  AND2X2 U1534 ( .A(n3198), .B(n7400), .Y(n7410) );
  AND2X2 U1535 ( .A(n3199), .B(n7410), .Y(n7420) );
  AND2X2 U1536 ( .A(n3200), .B(n7420), .Y(n7430) );
  AND2X2 U1537 ( .A(n3201), .B(n7430), .Y(n7440) );
  AND2X2 U1538 ( .A(n3202), .B(n7440), .Y(n7450) );
  AND2X2 U1539 ( .A(n3203), .B(n7450), .Y(n7460) );
  AND2X2 U1540 ( .A(n3204), .B(n7460), .Y(n7470) );
  AND2X2 U1541 ( .A(n3208), .B(n7370), .Y(n7480) );
  CLKINVX1 U1542 ( .A(stg4_real[16]), .Y(n1413) );
  CLKBUFX3 U1543 ( .A(n106), .Y(n853) );
  CLKBUFX3 U1544 ( .A(n106), .Y(n854) );
  CLKINVX1 U1545 ( .A(n1284), .Y(n1417) );
  AND2X2 U1546 ( .A(n3154), .B(n7610), .Y(n7490) );
  AND2X2 U1547 ( .A(n3185), .B(n7620), .Y(n7500) );
  AND2X2 U1548 ( .A(n3170), .B(n7630), .Y(n7510) );
  AND2X2 U1549 ( .A(n3156), .B(n7640), .Y(n7520) );
  AND2X2 U1550 ( .A(n3187), .B(n7650), .Y(n7530) );
  AND2X2 U1551 ( .A(n3172), .B(n7660), .Y(n7540) );
  CLKBUFX3 U1552 ( .A(n153), .Y(n911) );
  AND2X2 U1553 ( .A(n3151), .B(n3150), .Y(n7550) );
  AND2X2 U1554 ( .A(n3182), .B(n3181), .Y(n7560) );
  AND2X2 U1555 ( .A(n3167), .B(n3166), .Y(n7570) );
  AND2X2 U1556 ( .A(n3152), .B(n7550), .Y(n7580) );
  AND2X2 U1557 ( .A(n3183), .B(n7560), .Y(n7590) );
  AND2X2 U1558 ( .A(n3168), .B(n7570), .Y(n7600) );
  AND2X2 U1559 ( .A(n3153), .B(n7580), .Y(n7610) );
  AND2X2 U1560 ( .A(n3184), .B(n7590), .Y(n7620) );
  AND2X2 U1561 ( .A(n3169), .B(n7600), .Y(n7630) );
  AND2X2 U1562 ( .A(n3155), .B(n7490), .Y(n7640) );
  AND2X2 U1563 ( .A(n3186), .B(n7500), .Y(n7650) );
  AND2X2 U1564 ( .A(n3171), .B(n7510), .Y(n7660) );
  AND2X2 U1565 ( .A(n3157), .B(n7520), .Y(n7670) );
  AND2X2 U1566 ( .A(n3188), .B(n7530), .Y(n7680) );
  AND2X2 U1567 ( .A(n3173), .B(n7540), .Y(n7690) );
  AND2X2 U1568 ( .A(n3158), .B(n7670), .Y(n7700) );
  AND2X2 U1569 ( .A(n3189), .B(n7680), .Y(n7710) );
  AND2X2 U1570 ( .A(n3174), .B(n7690), .Y(n7720) );
  AND2X2 U1571 ( .A(n3159), .B(n7700), .Y(n7730) );
  AND2X2 U1572 ( .A(n3190), .B(n7710), .Y(n7740) );
  AND2X2 U1573 ( .A(n3175), .B(n7720), .Y(n7750) );
  AND2X2 U1574 ( .A(n3160), .B(n7730), .Y(n7760) );
  AND2X2 U1575 ( .A(n3191), .B(n7740), .Y(n7770) );
  AND2X2 U1576 ( .A(n3176), .B(n7750), .Y(n7780) );
  AND2X2 U1577 ( .A(n3161), .B(n7760), .Y(n7790) );
  AND2X2 U1578 ( .A(n3192), .B(n7770), .Y(n7800) );
  AND2X2 U1579 ( .A(n3177), .B(n7780), .Y(n7810) );
  AND2X2 U1580 ( .A(n3162), .B(n7790), .Y(n7820) );
  AND2X2 U1581 ( .A(n3193), .B(n7800), .Y(n7830) );
  AND2X2 U1582 ( .A(n3178), .B(n7810), .Y(n7840) );
  AND2X2 U1583 ( .A(n3163), .B(n7820), .Y(n7850) );
  AND2X2 U1584 ( .A(n2887), .B(n7830), .Y(n7860) );
  AND2X2 U1585 ( .A(n3179), .B(n7840), .Y(n7870) );
  CLKBUFX3 U1586 ( .A(n153), .Y(n910) );
  CLKBUFX3 U1587 ( .A(n2687), .Y(n851) );
  CLKBUFX3 U1588 ( .A(n7270), .Y(n9290) );
  AND2X2 U1589 ( .A(n3164), .B(n7850), .Y(n7880) );
  AND2X2 U1590 ( .A(n2876), .B(n7860), .Y(n7890) );
  AND2X2 U1591 ( .A(n3180), .B(n7870), .Y(n7900) );
  CLKBUFX3 U1592 ( .A(n7280), .Y(n868) );
  CLKBUFX3 U1593 ( .A(n7260), .Y(n912) );
  CLKBUFX3 U1594 ( .A(n7290), .Y(n9830) );
  OAI222XL U1595 ( .A0(n205), .A1(n2390), .B0(n850), .B1(n2870), .C0(n82), 
        .C1(n3081), .Y(n2020) );
  OAI222XL U1596 ( .A0(n195), .A1(n2394), .B0(n850), .B1(n2881), .C0(n83), 
        .C1(n2878), .Y(n2021) );
  OAI222XL U1597 ( .A0(n189), .A1(n2398), .B0(n850), .B1(n2893), .C0(n84), 
        .C1(n2889), .Y(n2022) );
  OAI222XL U1598 ( .A0(n181), .A1(n2402), .B0(n850), .B1(n2906), .C0(n80), 
        .C1(n2900), .Y(n2023) );
  OAI222XL U1599 ( .A0(n191), .A1(n2406), .B0(n849), .B1(n2919), .C0(n82), 
        .C1(n2913), .Y(n2024) );
  OAI222XL U1600 ( .A0(n193), .A1(n2410), .B0(n849), .B1(n2932), .C0(n81), 
        .C1(n2926), .Y(n2025) );
  OAI222XL U1601 ( .A0(n189), .A1(n2414), .B0(n849), .B1(n2945), .C0(n83), 
        .C1(n2939), .Y(n2026) );
  OAI222XL U1602 ( .A0(n3081), .A1(n864), .B0(n858), .B1(n2468), .C0(n205), 
        .C1(n2467), .Y(n1829) );
  OAI222XL U1603 ( .A0(n866), .A1(n2878), .B0(n858), .B1(n2473), .C0(n187), 
        .C1(n2472), .Y(n1830) );
  OAI222XL U1604 ( .A0(n865), .A1(n2889), .B0(n858), .B1(n2478), .C0(n189), 
        .C1(n2477), .Y(n1831) );
  OAI222XL U1605 ( .A0(n866), .A1(n2900), .B0(n858), .B1(n2483), .C0(n207), 
        .C1(n2482), .Y(n1832) );
  OAI222XL U1606 ( .A0(n866), .A1(n2913), .B0(n857), .B1(n2488), .C0(n197), 
        .C1(n2487), .Y(n1833) );
  OAI222XL U1607 ( .A0(n866), .A1(n2926), .B0(n857), .B1(n2493), .C0(n183), 
        .C1(n2492), .Y(n1834) );
  OAI222XL U1608 ( .A0(n865), .A1(n2939), .B0(n857), .B1(n2498), .C0(n200), 
        .C1(n2497), .Y(n1835) );
  OAI222XL U1609 ( .A0(n3081), .A1(n915), .B0(n911), .B1(n3084), .C0(n189), 
        .C1(n3083), .Y(n1924) );
  OAI222XL U1610 ( .A0(n912), .A1(n2878), .B0(n911), .B1(n3086), .C0(n193), 
        .C1(n2879), .Y(n1925) );
  OAI222XL U1611 ( .A0(n912), .A1(n2889), .B0(n911), .B1(n3088), .C0(n191), 
        .C1(n2890), .Y(n1926) );
  OAI222XL U1612 ( .A0(n912), .A1(n2900), .B0(n911), .B1(n3091), .C0(n202), 
        .C1(n2901), .Y(n1927) );
  OAI222XL U1613 ( .A0(n912), .A1(n2913), .B0(n910), .B1(n3095), .C0(n205), 
        .C1(n2914), .Y(n1928) );
  OAI222XL U1614 ( .A0(n912), .A1(n2926), .B0(n910), .B1(n3099), .C0(n183), 
        .C1(n2927), .Y(n1929) );
  OAI222XL U1615 ( .A0(n912), .A1(n2939), .B0(n910), .B1(n3103), .C0(n199), 
        .C1(n2940), .Y(n1930) );
  NAND4X2 U1616 ( .A(n3078), .B(n3077), .C(n3076), .D(n3075), .Y(mul_2_in[15])
         );
  OA22X1 U1617 ( .A0(n76), .A1(n3074), .B0(n10460), .B1(n3073), .Y(n3075) );
  OA22X1 U1618 ( .A0(n45), .A1(n91), .B0(n183), .B1(n96), .Y(n3076) );
  OA22X1 U1619 ( .A0(n9280), .A1(n89), .B0(n918), .B1(n90), .Y(n3077) );
  NAND4X2 U1620 ( .A(n2874), .B(n2873), .C(n2872), .D(n2871), .Y(mul_1_in[15])
         );
  OA22X1 U1621 ( .A0(n78), .A1(n2870), .B0(n10460), .B1(n2869), .Y(n2871) );
  OA22X1 U1622 ( .A0(n46), .A1(n113), .B0(n208), .B1(n2868), .Y(n2872) );
  OA22X1 U1623 ( .A0(n97), .A1(n9280), .B0(n917), .B1(n111), .Y(n2873) );
  OAI221XL U1624 ( .A0(n912), .A1(n3071), .B0(n200), .B1(n3070), .C0(n3069), 
        .Y(n1908) );
  AOI2BB2X1 U1625 ( .B0(stg2_real_6__15_), .B1(n869), .A0N(n911), .A1N(n3068), 
        .Y(n3069) );
  OAI221XL U1626 ( .A0(n915), .A1(n2711), .B0(n9690), .B1(n2710), .C0(n2709), 
        .Y(n1909) );
  AOI2BB2X1 U1627 ( .B0(stg2_real_6__14_), .B1(n875), .A0N(n911), .A1N(n2708), 
        .Y(n2709) );
  OAI221XL U1628 ( .A0(n912), .A1(n2573), .B0(n202), .B1(n1304), .C0(n1302), 
        .Y(n1910) );
  AOI2BB2X1 U1629 ( .B0(stg2_real_6__13_), .B1(n875), .A0N(n910), .A1N(n1306), 
        .Y(n1302) );
  OAI221XL U1630 ( .A0(n912), .A1(n2582), .B0(n202), .B1(n1313), .C0(n1311), 
        .Y(n1911) );
  AOI2BB2X1 U1631 ( .B0(stg2_real_6__12_), .B1(n876), .A0N(n910), .A1N(n1315), 
        .Y(n1311) );
  OAI221XL U1632 ( .A0(n912), .A1(n2591), .B0(n185), .B1(n1322), .C0(n1320), 
        .Y(n1912) );
  AOI2BB2X1 U1633 ( .B0(stg2_real_6__11_), .B1(n874), .A0N(n910), .A1N(n1324), 
        .Y(n1320) );
  OAI221XL U1634 ( .A0(n912), .A1(n2600), .B0(n187), .B1(n1331), .C0(n1329), 
        .Y(n1913) );
  AOI2BB2X1 U1635 ( .B0(stg2_real_6__10_), .B1(n874), .A0N(n910), .A1N(n1333), 
        .Y(n1329) );
  OAI221XL U1636 ( .A0(n912), .A1(n2609), .B0(n191), .B1(n1340), .C0(n1338), 
        .Y(n1914) );
  AOI2BB2X1 U1637 ( .B0(stg2_real_6__9_), .B1(n874), .A0N(n910), .A1N(n1342), 
        .Y(n1338) );
  OAI221XL U1638 ( .A0(n864), .A1(n3071), .B0(n203), .B1(n2558), .C0(n2556), 
        .Y(n1813) );
  AOI2BB2X1 U1639 ( .B0(stg2_real_7__15_), .B1(n873), .A0N(n858), .A1N(n2560), 
        .Y(n2556) );
  OAI221XL U1640 ( .A0(n864), .A1(n2711), .B0(n202), .B1(n2566), .C0(n2564), 
        .Y(n1814) );
  AOI2BB2X1 U1641 ( .B0(stg2_real_7__14_), .B1(n875), .A0N(n858), .A1N(n2568), 
        .Y(n2564) );
  OAI221XL U1642 ( .A0(n864), .A1(n2573), .B0(n205), .B1(n2575), .C0(n2572), 
        .Y(n1815) );
  AOI2BB2X1 U1643 ( .B0(stg2_real_7__13_), .B1(n874), .A0N(n858), .A1N(n2577), 
        .Y(n2572) );
  OAI221XL U1644 ( .A0(n864), .A1(n2582), .B0(n207), .B1(n2584), .C0(n2581), 
        .Y(n1816) );
  AOI2BB2X1 U1645 ( .B0(stg2_real_7__12_), .B1(n874), .A0N(n858), .A1N(n2586), 
        .Y(n2581) );
  OAI221XL U1646 ( .A0(n865), .A1(n2591), .B0(n183), .B1(n2593), .C0(n2590), 
        .Y(n1817) );
  AOI2BB2X1 U1647 ( .B0(stg2_real_7__11_), .B1(n874), .A0N(n858), .A1N(n2595), 
        .Y(n2590) );
  OAI221XL U1648 ( .A0(n864), .A1(n2600), .B0(n181), .B1(n2602), .C0(n2599), 
        .Y(n1818) );
  AOI2BB2X1 U1649 ( .B0(stg2_real_7__10_), .B1(n872), .A0N(n857), .A1N(n2604), 
        .Y(n2599) );
  OAI221XL U1650 ( .A0(n865), .A1(n2609), .B0(n197), .B1(n2611), .C0(n2608), 
        .Y(n1819) );
  AOI2BB2X1 U1651 ( .B0(stg2_real_7__9_), .B1(n875), .A0N(n858), .A1N(n2613), 
        .Y(n2608) );
  AOI2BB2X1 U1652 ( .B0(stg2_img_15__15_), .B1(n873), .A0N(n3081), .A1N(n852), 
        .Y(n2464) );
  OAI221XL U1653 ( .A0(n9290), .A1(n2472), .B0(n854), .B1(n2880), .C0(n2470), 
        .Y(n1862) );
  AOI2BB2X1 U1654 ( .B0(stg2_img_15__14_), .B1(n873), .A0N(n2878), .A1N(n851), 
        .Y(n2470) );
  XOR2X1 U1655 ( .A(n3208), .B(n7370), .Y(stg2_img_15__14_) );
  OAI221XL U1656 ( .A0(n9290), .A1(n2477), .B0(n854), .B1(n2892), .C0(n2475), 
        .Y(n1863) );
  XOR2X1 U1657 ( .A(n3207), .B(n7360), .Y(stg2_img_15__13_) );
  OAI221XL U1658 ( .A0(n9340), .A1(n2482), .B0(n854), .B1(n2905), .C0(n2480), 
        .Y(n1864) );
  XOR2X1 U1659 ( .A(n3206), .B(n7350), .Y(stg2_img_15__12_) );
  OAI221XL U1660 ( .A0(n9330), .A1(n2487), .B0(n854), .B1(n2918), .C0(n2485), 
        .Y(n1865) );
  XOR2X1 U1661 ( .A(n3205), .B(n7470), .Y(stg2_img_15__11_) );
  OAI221XL U1662 ( .A0(n9290), .A1(n2492), .B0(n854), .B1(n2931), .C0(n2490), 
        .Y(n1866) );
  XOR2X1 U1663 ( .A(n3204), .B(n7460), .Y(stg2_img_15__10_) );
  OAI221XL U1664 ( .A0(n9290), .A1(n2497), .B0(n854), .B1(n2944), .C0(n2495), 
        .Y(n1867) );
  XOR2X1 U1665 ( .A(n3203), .B(n7450), .Y(stg2_img_15__9_) );
  OAI221XL U1666 ( .A0(n9290), .A1(n2502), .B0(n854), .B1(n2957), .C0(n2500), 
        .Y(n1868) );
  XOR2X1 U1667 ( .A(n3202), .B(n7440), .Y(stg2_img_15__8_) );
  OAI221XL U1668 ( .A0(n9330), .A1(n2575), .B0(n853), .B1(n2725), .C0(n2570), 
        .Y(n1847) );
  OAI221XL U1669 ( .A0(n9330), .A1(n2584), .B0(n106), .B1(n2735), .C0(n2579), 
        .Y(n1848) );
  OAI221XL U1670 ( .A0(n9340), .A1(n2593), .B0(n853), .B1(n2745), .C0(n2588), 
        .Y(n1849) );
  OAI221XL U1671 ( .A0(n9340), .A1(n2602), .B0(n853), .B1(n2755), .C0(n2597), 
        .Y(n1850) );
  OAI221XL U1672 ( .A0(n9330), .A1(n2611), .B0(n853), .B1(n2765), .C0(n2606), 
        .Y(n1851) );
  OAI221XL U1673 ( .A0(n9330), .A1(n2620), .B0(n853), .B1(n2775), .C0(n2615), 
        .Y(n1852) );
  OAI221XL U1674 ( .A0(n9340), .A1(n2629), .B0(n853), .B1(n2785), .C0(n2624), 
        .Y(n1853) );
  AOI2BB2X1 U1675 ( .B0(stg2_real_5__15_), .B1(n872), .A0N(n850), .A1N(n3074), 
        .Y(n1423) );
  OAI221XL U1676 ( .A0(n203), .A1(n1432), .B0(n80), .B1(n2711), .C0(n1430), 
        .Y(n2005) );
  AOI2BB2X1 U1677 ( .B0(stg2_real_5__14_), .B1(n872), .A0N(n849), .A1N(n2716), 
        .Y(n1430) );
  OAI221XL U1678 ( .A0(n207), .A1(n1795), .B0(n79), .B1(n2573), .C0(n1793), 
        .Y(n2006) );
  AOI2BB2X1 U1679 ( .B0(stg2_real_5__13_), .B1(n872), .A0N(n849), .A1N(n2726), 
        .Y(n1793) );
  OAI221XL U1680 ( .A0(n197), .A1(n1802), .B0(n78), .B1(n2582), .C0(n1800), 
        .Y(n2007) );
  AOI2BB2X1 U1681 ( .B0(stg2_real_5__12_), .B1(n873), .A0N(n849), .A1N(n2736), 
        .Y(n1800) );
  OAI221XL U1682 ( .A0(n205), .A1(n1809), .B0(n79), .B1(n2591), .C0(n1807), 
        .Y(n2008) );
  AOI2BB2X1 U1683 ( .B0(stg2_real_5__11_), .B1(n871), .A0N(n849), .A1N(n2746), 
        .Y(n1807) );
  OAI221XL U1684 ( .A0(n189), .A1(n2314), .B0(n78), .B1(n2600), .C0(n2312), 
        .Y(n2009) );
  AOI2BB2X1 U1685 ( .B0(stg2_real_5__10_), .B1(n871), .A0N(n849), .A1N(n2756), 
        .Y(n2312) );
  OAI221XL U1686 ( .A0(n195), .A1(n2321), .B0(n81), .B1(n2609), .C0(n2319), 
        .Y(n2010) );
  AOI2BB2X1 U1687 ( .B0(stg2_real_5__9_), .B1(n871), .A0N(n849), .A1N(n2766), 
        .Y(n2319) );
  OAI221XL U1688 ( .A0(n185), .A1(n2328), .B0(n77), .B1(n2618), .C0(n2326), 
        .Y(n2011) );
  AOI2BB2X1 U1689 ( .B0(stg2_real_5__8_), .B1(n871), .A0N(n850), .A1N(n2776), 
        .Y(n2326) );
  OAI221XL U1690 ( .A0(n909), .A1(n3071), .B0(n52), .B1(n3070), .C0(n1288), 
        .Y(n1972) );
  AOI2BB1X1 U1691 ( .A0N(n902), .A1N(n152), .B0(n103), .Y(n1288) );
  OAI221XL U1692 ( .A0(n909), .A1(n2711), .B0(n20), .B1(n2710), .C0(n1293), 
        .Y(n1973) );
  AOI2BB1X1 U1693 ( .A0N(n901), .A1N(n1297), .B0(n808), .Y(n1293) );
  OAI221XL U1694 ( .A0(n909), .A1(n2573), .B0(n48), .B1(n1304), .C0(n1299), 
        .Y(n1974) );
  AOI2BB1X1 U1695 ( .A0N(n901), .A1N(n1308), .B0(n809), .Y(n1299) );
  OAI221XL U1696 ( .A0(n908), .A1(n2582), .B0(n47), .B1(n1313), .C0(n1310), 
        .Y(n1975) );
  AOI2BB1X1 U1697 ( .A0N(n901), .A1N(n1317), .B0(n810), .Y(n1310) );
  OAI221XL U1698 ( .A0(n908), .A1(n2591), .B0(n51), .B1(n1322), .C0(n1319), 
        .Y(n1976) );
  AOI2BB1X1 U1699 ( .A0N(n901), .A1N(n1326), .B0(n811), .Y(n1319) );
  OAI221XL U1700 ( .A0(n908), .A1(n2600), .B0(n49), .B1(n1331), .C0(n1328), 
        .Y(n1977) );
  AOI2BB1X1 U1701 ( .A0N(n901), .A1N(n1335), .B0(n812), .Y(n1328) );
  OAI221XL U1702 ( .A0(n908), .A1(n2609), .B0(n45), .B1(n1340), .C0(n1337), 
        .Y(n1978) );
  AOI2BB1X1 U1703 ( .A0N(n902), .A1N(n1344), .B0(n813), .Y(n1337) );
  OAI221XL U1704 ( .A0(n917), .A1(n3071), .B0(n48), .B1(n2558), .C0(n2555), 
        .Y(n1876) );
  AOI2BB1X1 U1705 ( .A0N(n855), .A1N(n90), .B0(n104), .Y(n2555) );
  OAI221XL U1706 ( .A0(n917), .A1(n2711), .B0(n47), .B1(n2566), .C0(n2563), 
        .Y(n1877) );
  AOI2BB1X1 U1707 ( .A0N(n855), .A1N(n2712), .B0(n822), .Y(n2563) );
  OAI221XL U1708 ( .A0(n9200), .A1(n2573), .B0(n50), .B1(n2575), .C0(n2571), 
        .Y(n1878) );
  AOI2BB1X1 U1709 ( .A0N(n855), .A1N(n2721), .B0(n832), .Y(n2571) );
  OAI221XL U1710 ( .A0(n917), .A1(n2582), .B0(n50), .B1(n2584), .C0(n2580), 
        .Y(n1879) );
  AOI2BB1X1 U1711 ( .A0N(n855), .A1N(n2731), .B0(n833), .Y(n2580) );
  OAI221XL U1712 ( .A0(n917), .A1(n2591), .B0(n48), .B1(n2593), .C0(n2589), 
        .Y(n1880) );
  AOI2BB1X1 U1713 ( .A0N(n855), .A1N(n2741), .B0(n834), .Y(n2589) );
  OAI221XL U1714 ( .A0(n917), .A1(n2600), .B0(n51), .B1(n2602), .C0(n2598), 
        .Y(n1881) );
  AOI2BB1X1 U1715 ( .A0N(n855), .A1N(n2751), .B0(n823), .Y(n2598) );
  OAI221XL U1716 ( .A0(n917), .A1(n2609), .B0(n49), .B1(n2611), .C0(n2607), 
        .Y(n1882) );
  AOI2BB1X1 U1717 ( .A0N(n856), .A1N(n2761), .B0(n824), .Y(n2607) );
  OAI221XL U1718 ( .A0(n3083), .A1(n9310), .B0(n9270), .B1(n3081), .C0(n3080), 
        .Y(n1956) );
  AOI2BB2X1 U1719 ( .B0(stg2_img_14__15_), .B1(n874), .A0N(n9230), .A1N(n97), 
        .Y(n3080) );
  OAI221XL U1720 ( .A0(n2879), .A1(n9300), .B0(n9270), .B1(n2878), .C0(n2877), 
        .Y(n1957) );
  AOI2BB2X1 U1721 ( .B0(stg2_img_14__14_), .B1(n869), .A0N(n9230), .A1N(n94), 
        .Y(n2877) );
  XOR2X1 U1722 ( .A(n2876), .B(n7860), .Y(stg2_img_14__14_) );
  OAI221XL U1723 ( .A0(n2890), .A1(n9290), .B0(n9270), .B1(n2889), .C0(n2888), 
        .Y(n1958) );
  AOI2BB2X1 U1724 ( .B0(stg2_img_14__13_), .B1(n876), .A0N(n9240), .A1N(n3090), 
        .Y(n2888) );
  XOR2X1 U1725 ( .A(n2887), .B(n7830), .Y(stg2_img_14__13_) );
  OAI221XL U1726 ( .A0(n2901), .A1(n9300), .B0(n9270), .B1(n2900), .C0(n2899), 
        .Y(n1959) );
  AOI2BB2X1 U1727 ( .B0(stg2_img_14__12_), .B1(n869), .A0N(n9240), .A1N(n3094), 
        .Y(n2899) );
  XOR2X1 U1728 ( .A(n3193), .B(n7800), .Y(stg2_img_14__12_) );
  OAI221XL U1729 ( .A0(n2914), .A1(n9300), .B0(n9270), .B1(n2913), .C0(n2912), 
        .Y(n1960) );
  AOI2BB2X1 U1730 ( .B0(stg2_img_14__11_), .B1(n869), .A0N(n9230), .A1N(n3098), 
        .Y(n2912) );
  XOR2X1 U1731 ( .A(n3192), .B(n7770), .Y(stg2_img_14__11_) );
  OAI221XL U1732 ( .A0(n2927), .A1(n9300), .B0(n9270), .B1(n2926), .C0(n2925), 
        .Y(n1961) );
  AOI2BB2X1 U1733 ( .B0(stg2_img_14__10_), .B1(n874), .A0N(n9240), .A1N(n3102), 
        .Y(n2925) );
  XOR2X1 U1734 ( .A(n3191), .B(n7740), .Y(stg2_img_14__10_) );
  OAI221XL U1735 ( .A0(n2940), .A1(n9350), .B0(n9270), .B1(n2939), .C0(n2938), 
        .Y(n1962) );
  AOI2BB2X1 U1736 ( .B0(stg2_img_14__9_), .B1(n869), .A0N(n9230), .A1N(n3106), 
        .Y(n2938) );
  XOR2X1 U1737 ( .A(n3190), .B(n7710), .Y(stg2_img_14__9_) );
  AOI2BB1X1 U1738 ( .A0N(n848), .A1N(n96), .B0(n120), .Y(n1422) );
  OAI221XL U1739 ( .A0(n9350), .A1(n2710), .B0(n9260), .B1(n2711), .C0(n1292), 
        .Y(n1941) );
  AOI2BB1X1 U1740 ( .A0N(n9240), .A1N(n2713), .B0(n808), .Y(n1292) );
  OAI221XL U1741 ( .A0(n9350), .A1(n1304), .B0(n9260), .B1(n2573), .C0(n1298), 
        .Y(n1942) );
  AOI2BB1X1 U1742 ( .A0N(n9230), .A1N(n2722), .B0(n809), .Y(n1298) );
  OAI221XL U1743 ( .A0(n9350), .A1(n1313), .B0(n9260), .B1(n2582), .C0(n1309), 
        .Y(n1943) );
  AOI2BB1X1 U1744 ( .A0N(n9240), .A1N(n2732), .B0(n810), .Y(n1309) );
  OAI221XL U1745 ( .A0(n9350), .A1(n1322), .B0(n9260), .B1(n2591), .C0(n1318), 
        .Y(n1944) );
  AOI2BB1X1 U1746 ( .A0N(n9230), .A1N(n2742), .B0(n811), .Y(n1318) );
  OAI221XL U1747 ( .A0(n9350), .A1(n1331), .B0(n9260), .B1(n2600), .C0(n1327), 
        .Y(n1945) );
  AOI2BB1X1 U1748 ( .A0N(n3079), .A1N(n2752), .B0(n812), .Y(n1327) );
  OAI221XL U1749 ( .A0(n9320), .A1(n1340), .B0(n9260), .B1(n2609), .C0(n1336), 
        .Y(n1946) );
  AOI2BB1X1 U1750 ( .A0N(n3079), .A1N(n2762), .B0(n813), .Y(n1336) );
  AOI2BB1X1 U1751 ( .A0N(n846), .A1N(n91), .B0(n120), .Y(n1419) );
  OAI221XL U1752 ( .A0(n52), .A1(n1432), .B0(n193), .B1(n2711), .C0(n1429), 
        .Y(n2069) );
  AOI2BB1X1 U1753 ( .A0N(n847), .A1N(n92), .B0(n794), .Y(n1429) );
  AOI2BB1X1 U1754 ( .A0N(n9240), .A1N(n89), .B0(n103), .Y(n1286) );
  OAI221XL U1755 ( .A0(n9300), .A1(n1432), .B0(n51), .B1(n2711), .C0(n1428), 
        .Y(n2037) );
  AOI2BB1X1 U1756 ( .A0N(n2456), .A1N(n2714), .B0(n794), .Y(n1428) );
  OAI221XL U1757 ( .A0(n20), .A1(n1795), .B0(n195), .B1(n2573), .C0(n1436), 
        .Y(n2070) );
  AOI2BB1X1 U1758 ( .A0N(n847), .A1N(n2723), .B0(n795), .Y(n1436) );
  OAI221XL U1759 ( .A0(n9320), .A1(n1795), .B0(n46), .B1(n2573), .C0(n1435), 
        .Y(n2038) );
  AOI2BB1X1 U1760 ( .A0N(n845), .A1N(n2724), .B0(n795), .Y(n1435) );
  OAI221XL U1761 ( .A0(n45), .A1(n1802), .B0(n200), .B1(n2582), .C0(n1799), 
        .Y(n2071) );
  AOI2BB1X1 U1762 ( .A0N(n847), .A1N(n2733), .B0(n796), .Y(n1799) );
  OAI221XL U1763 ( .A0(n9310), .A1(n1802), .B0(n20), .B1(n2582), .C0(n1798), 
        .Y(n2039) );
  AOI2BB1X1 U1764 ( .A0N(n846), .A1N(n2734), .B0(n796), .Y(n1798) );
  OAI221XL U1765 ( .A0(n19), .A1(n1809), .B0(n195), .B1(n2591), .C0(n1806), 
        .Y(n2072) );
  AOI2BB1X1 U1766 ( .A0N(n847), .A1N(n2743), .B0(n797), .Y(n1806) );
  OAI221XL U1767 ( .A0(n9320), .A1(n1809), .B0(n51), .B1(n2591), .C0(n1805), 
        .Y(n2040) );
  AOI2BB1X1 U1768 ( .A0N(n845), .A1N(n2744), .B0(n797), .Y(n1805) );
  OAI221XL U1769 ( .A0(n19), .A1(n2314), .B0(n199), .B1(n2600), .C0(n2311), 
        .Y(n2073) );
  AOI2BB1X1 U1770 ( .A0N(n847), .A1N(n2753), .B0(n798), .Y(n2311) );
  OAI221XL U1771 ( .A0(n9290), .A1(n2314), .B0(n47), .B1(n2600), .C0(n2310), 
        .Y(n2041) );
  AOI2BB1X1 U1772 ( .A0N(n2456), .A1N(n2754), .B0(n798), .Y(n2310) );
  OAI221XL U1773 ( .A0(n20), .A1(n2321), .B0(n189), .B1(n2609), .C0(n2318), 
        .Y(n2074) );
  AOI2BB1X1 U1774 ( .A0N(n848), .A1N(n2763), .B0(n799), .Y(n2318) );
  OAI221XL U1775 ( .A0(n9310), .A1(n2321), .B0(n19), .B1(n2609), .C0(n2317), 
        .Y(n2042) );
  AOI2BB1X1 U1776 ( .A0N(n2456), .A1N(n2764), .B0(n799), .Y(n2317) );
  OAI221XL U1777 ( .A0(n9290), .A1(n2390), .B0(n52), .B1(n3081), .C0(n2387), 
        .Y(n2052) );
  AOI2BB2X1 U1778 ( .B0(stg2_img_13__15_), .B1(n870), .A0N(n846), .A1N(n113), 
        .Y(n2387) );
  OAI221XL U1779 ( .A0(n9320), .A1(n2394), .B0(n45), .B1(n2878), .C0(n2392), 
        .Y(n2053) );
  AOI2BB2X1 U1780 ( .B0(stg2_img_13__14_), .B1(n870), .A0N(n846), .A1N(n110), 
        .Y(n2392) );
  XOR2X1 U1781 ( .A(n3180), .B(n7870), .Y(stg2_img_13__14_) );
  OAI221XL U1782 ( .A0(n9310), .A1(n2398), .B0(n46), .B1(n2889), .C0(n2396), 
        .Y(n2054) );
  AOI2BB2X1 U1783 ( .B0(stg2_img_13__13_), .B1(n870), .A0N(n846), .A1N(n2891), 
        .Y(n2396) );
  XOR2X1 U1784 ( .A(n3179), .B(n7840), .Y(stg2_img_13__13_) );
  OAI221XL U1785 ( .A0(n9320), .A1(n2402), .B0(n47), .B1(n2900), .C0(n2400), 
        .Y(n2055) );
  AOI2BB2X1 U1786 ( .B0(stg2_img_13__12_), .B1(n870), .A0N(n845), .A1N(n2904), 
        .Y(n2400) );
  XOR2X1 U1787 ( .A(n3178), .B(n7810), .Y(stg2_img_13__12_) );
  OAI221XL U1788 ( .A0(n9290), .A1(n2406), .B0(n19), .B1(n2913), .C0(n2404), 
        .Y(n2056) );
  AOI2BB2X1 U1789 ( .B0(stg2_img_13__11_), .B1(n870), .A0N(n845), .A1N(n2917), 
        .Y(n2404) );
  XOR2X1 U1790 ( .A(n3177), .B(n7780), .Y(stg2_img_13__11_) );
  OAI221XL U1791 ( .A0(n9320), .A1(n2410), .B0(n46), .B1(n2926), .C0(n2408), 
        .Y(n2057) );
  AOI2BB2X1 U1792 ( .B0(stg2_img_13__10_), .B1(n870), .A0N(n845), .A1N(n2930), 
        .Y(n2408) );
  XOR2X1 U1793 ( .A(n3176), .B(n7750), .Y(stg2_img_13__10_) );
  OAI221XL U1794 ( .A0(n9320), .A1(n2414), .B0(n49), .B1(n2939), .C0(n2412), 
        .Y(n2058) );
  AOI2BB2X1 U1795 ( .B0(stg2_img_13__9_), .B1(n870), .A0N(n845), .A1N(n2943), 
        .Y(n2412) );
  XOR2X1 U1796 ( .A(n3175), .B(n7720), .Y(stg2_img_13__9_) );
  CLKINVX1 U1797 ( .A(stg2_img_11__15_), .Y(n2466) );
  OA22X1 U1798 ( .A0(n3081), .A1(n917), .B0(n45), .B1(n2467), .Y(n2465) );
  OAI221XL U1799 ( .A0(n855), .A1(n112), .B0(n893), .B1(n3208), .C0(n2471), 
        .Y(n1893) );
  OA22X1 U1800 ( .A0(n917), .A1(n2878), .B0(n45), .B1(n2472), .Y(n2471) );
  OAI221XL U1801 ( .A0(n855), .A1(n108), .B0(n893), .B1(n3207), .C0(n2476), 
        .Y(n1894) );
  OA22X1 U1802 ( .A0(n9190), .A1(n2889), .B0(n47), .B1(n2477), .Y(n2476) );
  OAI221XL U1803 ( .A0(n855), .A1(n2902), .B0(n892), .B1(n3206), .C0(n2481), 
        .Y(n1895) );
  OAI221XL U1804 ( .A0(n855), .A1(n2915), .B0(n892), .B1(n3205), .C0(n2486), 
        .Y(n1896) );
  OAI221XL U1805 ( .A0(n855), .A1(n2928), .B0(n892), .B1(n3204), .C0(n2491), 
        .Y(n1897) );
  OAI221XL U1806 ( .A0(n855), .A1(n2941), .B0(n892), .B1(n3203), .C0(n2496), 
        .Y(n1898) );
  OAI221XL U1807 ( .A0(n855), .A1(n2954), .B0(n892), .B1(n3202), .C0(n2501), 
        .Y(n1899) );
  OAI221XL U1808 ( .A0(n901), .A1(n3093), .B0(n890), .B1(n3193), .C0(n2898), 
        .Y(n1991) );
  OAI221XL U1809 ( .A0(n901), .A1(n3110), .B0(n889), .B1(n3189), .C0(n2950), 
        .Y(n1995) );
  CLKINVX1 U1810 ( .A(stg2_img_9__15_), .Y(n2389) );
  OA22X1 U1811 ( .A0(n49), .A1(n2390), .B0(n189), .B1(n3081), .Y(n2388) );
  OAI221XL U1812 ( .A0(n848), .A1(n95), .B0(n895), .B1(n3180), .C0(n2393), .Y(
        n2085) );
  OA22X1 U1813 ( .A0(n48), .A1(n2394), .B0(n199), .B1(n2878), .Y(n2393) );
  OAI221XL U1814 ( .A0(n848), .A1(n93), .B0(n895), .B1(n3179), .C0(n2397), .Y(
        n2086) );
  OAI221XL U1815 ( .A0(n847), .A1(n2903), .B0(n895), .B1(n3178), .C0(n2401), 
        .Y(n2087) );
  OAI221XL U1816 ( .A0(n847), .A1(n2916), .B0(n895), .B1(n3177), .C0(n2405), 
        .Y(n2088) );
  OAI221XL U1817 ( .A0(n847), .A1(n2929), .B0(n895), .B1(n3176), .C0(n2409), 
        .Y(n2089) );
  OAI221XL U1818 ( .A0(n847), .A1(n2942), .B0(n895), .B1(n3175), .C0(n2413), 
        .Y(n2090) );
  OAI221XL U1819 ( .A0(n847), .A1(n2955), .B0(n894), .B1(n3174), .C0(n2417), 
        .Y(n2091) );
  CLKINVX1 U1820 ( .A(n10500), .Y(n10480) );
  AND2X2 U1821 ( .A(n838), .B(n109), .Y(n791) );
  CLKINVX1 U1822 ( .A(stg2_img_10__15_), .Y(n2867) );
  OA22X1 U1823 ( .A0(n3081), .A1(n906), .B0(n46), .B1(n3083), .Y(n2866) );
  OAI221XL U1824 ( .A0(n902), .A1(n151), .B0(n891), .B1(n2876), .C0(n2875), 
        .Y(n1989) );
  CLKINVX1 U1825 ( .A(stg2_img_10__14_), .Y(n2876) );
  OA22X1 U1826 ( .A0(n909), .A1(n2878), .B0(n48), .B1(n2879), .Y(n2875) );
  OAI221XL U1827 ( .A0(n902), .A1(n132), .B0(n890), .B1(n2887), .C0(n2886), 
        .Y(n1990) );
  CLKINVX1 U1828 ( .A(stg2_img_10__13_), .Y(n2887) );
  OA22X1 U1829 ( .A0(n906), .A1(n2889), .B0(n48), .B1(n2890), .Y(n2886) );
  OAI221XL U1830 ( .A0(n901), .A1(n3097), .B0(n889), .B1(n3192), .C0(n2911), 
        .Y(n1992) );
  OAI221XL U1831 ( .A0(n901), .A1(n3101), .B0(n889), .B1(n3191), .C0(n2924), 
        .Y(n1993) );
  OAI221XL U1832 ( .A0(n901), .A1(n3105), .B0(n890), .B1(n3190), .C0(n2937), 
        .Y(n1994) );
  OA22X1 U1833 ( .A0(n202), .A1(n2696), .B0(n78), .B1(n2695), .Y(n2697) );
  OA22X1 U1834 ( .A0(n200), .A1(n2856), .B0(n75), .B1(n2385), .Y(n2386) );
  OAI222XL U1835 ( .A0(n199), .A1(n2418), .B0(n849), .B1(n2958), .C0(n81), 
        .C1(n2952), .Y(n2027) );
  OAI222XL U1836 ( .A0(n181), .A1(n2423), .B0(n849), .B1(n2971), .C0(n75), 
        .C1(n2965), .Y(n2028) );
  OAI222XL U1837 ( .A0(n191), .A1(n2428), .B0(n849), .B1(n2984), .C0(n84), 
        .C1(n2978), .Y(n2029) );
  OAI222XL U1838 ( .A0(n193), .A1(n2433), .B0(n849), .B1(n2997), .C0(n83), 
        .C1(n2991), .Y(n2030) );
  OAI222XL U1839 ( .A0(n199), .A1(n2438), .B0(n849), .B1(n3010), .C0(n80), 
        .C1(n3004), .Y(n2031) );
  OAI222XL U1840 ( .A0(n195), .A1(n2443), .B0(n849), .B1(n3023), .C0(n79), 
        .C1(n3017), .Y(n2032) );
  OAI222XL U1841 ( .A0(n187), .A1(n2448), .B0(n849), .B1(n3036), .C0(n77), 
        .C1(n3030), .Y(n2033) );
  OAI222XL U1842 ( .A0(n197), .A1(n2453), .B0(n849), .B1(n3049), .C0(n78), 
        .C1(n3043), .Y(n2034) );
  OAI222XL U1843 ( .A0(n181), .A1(n2461), .B0(n849), .B1(n3063), .C0(n76), 
        .C1(n3057), .Y(n2035) );
  OAI222XL U1844 ( .A0(n865), .A1(n2952), .B0(n857), .B1(n2504), .C0(n203), 
        .C1(n2502), .Y(n1836) );
  OAI222XL U1845 ( .A0(n865), .A1(n2965), .B0(n857), .B1(n2510), .C0(n207), 
        .C1(n2508), .Y(n1837) );
  OAI222XL U1846 ( .A0(n865), .A1(n2978), .B0(n857), .B1(n2516), .C0(n195), 
        .C1(n2514), .Y(n1838) );
  OAI222XL U1847 ( .A0(n865), .A1(n2991), .B0(n857), .B1(n2522), .C0(n197), 
        .C1(n2520), .Y(n1839) );
  OAI222XL U1848 ( .A0(n865), .A1(n3004), .B0(n857), .B1(n2528), .C0(n183), 
        .C1(n2526), .Y(n1840) );
  OAI222XL U1849 ( .A0(n865), .A1(n3017), .B0(n857), .B1(n2534), .C0(n187), 
        .C1(n2532), .Y(n1841) );
  OAI222XL U1850 ( .A0(n865), .A1(n3030), .B0(n857), .B1(n2540), .C0(n195), 
        .C1(n2538), .Y(n1842) );
  OAI222XL U1851 ( .A0(n864), .A1(n3043), .B0(n857), .B1(n2546), .C0(n199), 
        .C1(n2544), .Y(n1843) );
  OAI222XL U1852 ( .A0(n864), .A1(n3057), .B0(n857), .B1(n2552), .C0(n199), 
        .C1(n2550), .Y(n1844) );
  OAI222XL U1853 ( .A0(n912), .A1(n2952), .B0(n910), .B1(n3108), .C0(n185), 
        .C1(n2953), .Y(n1931) );
  OAI222XL U1854 ( .A0(n912), .A1(n2965), .B0(n910), .B1(n3113), .C0(n207), 
        .C1(n2966), .Y(n1932) );
  OAI222XL U1855 ( .A0(n912), .A1(n2978), .B0(n910), .B1(n3117), .C0(n181), 
        .C1(n2979), .Y(n1933) );
  OAI222XL U1856 ( .A0(n912), .A1(n2991), .B0(n910), .B1(n3122), .C0(n9650), 
        .C1(n2992), .Y(n1934) );
  OAI222XL U1857 ( .A0(n915), .A1(n3004), .B0(n910), .B1(n3127), .C0(n185), 
        .C1(n3005), .Y(n1935) );
  OAI222XL U1858 ( .A0(n915), .A1(n3017), .B0(n910), .B1(n3131), .C0(n187), 
        .C1(n3018), .Y(n1936) );
  OAI222XL U1859 ( .A0(n915), .A1(n3030), .B0(n910), .B1(n3135), .C0(n181), 
        .C1(n3031), .Y(n1937) );
  OAI222XL U1860 ( .A0(n915), .A1(n3043), .B0(n910), .B1(n3139), .C0(n191), 
        .C1(n3044), .Y(n1938) );
  OAI222XL U1861 ( .A0(n915), .A1(n3057), .B0(n910), .B1(n3145), .C0(n193), 
        .C1(n3058), .Y(n1939) );
  OAI221XL U1862 ( .A0(n915), .A1(n2692), .B0(n193), .B1(n1413), .C0(n1411), 
        .Y(n1923) );
  AOI2BB2X1 U1863 ( .B0(stg2_real_6__0_), .B1(n874), .A0N(n911), .A1N(n1415), 
        .Y(n1411) );
  OAI221XL U1864 ( .A0(n864), .A1(n2692), .B0(n203), .B1(n2694), .C0(n2691), 
        .Y(n1828) );
  AOI2BB2X1 U1865 ( .B0(stg2_real_7__0_), .B1(n869), .A0N(n858), .A1N(n2696), 
        .Y(n2691) );
  OAI221XL U1866 ( .A0(n912), .A1(n2618), .B0(n189), .B1(n1349), .C0(n1347), 
        .Y(n1915) );
  AOI2BB2X1 U1867 ( .B0(stg2_real_6__8_), .B1(n874), .A0N(n911), .A1N(n1351), 
        .Y(n1347) );
  OAI221XL U1868 ( .A0(n912), .A1(n2627), .B0(n185), .B1(n1357), .C0(n1355), 
        .Y(n1916) );
  AOI2BB2X1 U1869 ( .B0(stg2_real_6__7_), .B1(n875), .A0N(n911), .A1N(n1359), 
        .Y(n1355) );
  OAI221XL U1870 ( .A0(n915), .A1(n2636), .B0(n191), .B1(n1365), .C0(n1363), 
        .Y(n1917) );
  AOI2BB2X1 U1871 ( .B0(stg2_real_6__6_), .B1(n875), .A0N(n911), .A1N(n1367), 
        .Y(n1363) );
  OAI221XL U1872 ( .A0(n912), .A1(n2645), .B0(n199), .B1(n1373), .C0(n1371), 
        .Y(n1918) );
  AOI2BB2X1 U1873 ( .B0(stg2_real_6__5_), .B1(n873), .A0N(n911), .A1N(n1375), 
        .Y(n1371) );
  OAI221XL U1874 ( .A0(n912), .A1(n2654), .B0(n189), .B1(n1381), .C0(n1379), 
        .Y(n1919) );
  AOI2BB2X1 U1875 ( .B0(stg2_real_6__4_), .B1(n873), .A0N(n911), .A1N(n1383), 
        .Y(n1379) );
  OAI221XL U1876 ( .A0(n916), .A1(n2663), .B0(n187), .B1(n1389), .C0(n1387), 
        .Y(n1920) );
  AOI2BB2X1 U1877 ( .B0(stg2_real_6__3_), .B1(n873), .A0N(n911), .A1N(n1391), 
        .Y(n1387) );
  OAI221XL U1878 ( .A0(n916), .A1(n2672), .B0(n207), .B1(n1397), .C0(n1395), 
        .Y(n1921) );
  AOI2BB2X1 U1879 ( .B0(stg2_real_6__2_), .B1(n873), .A0N(n911), .A1N(n1399), 
        .Y(n1395) );
  OAI221XL U1880 ( .A0(n915), .A1(n2681), .B0(n181), .B1(n1405), .C0(n1403), 
        .Y(n1922) );
  AOI2BB2X1 U1881 ( .B0(stg2_real_6__1_), .B1(n873), .A0N(n911), .A1N(n1407), 
        .Y(n1403) );
  OAI221XL U1882 ( .A0(n864), .A1(n2618), .B0(n200), .B1(n2620), .C0(n2617), 
        .Y(n1820) );
  AOI2BB2X1 U1883 ( .B0(stg2_real_7__8_), .B1(n875), .A0N(n858), .A1N(n2622), 
        .Y(n2617) );
  OAI221XL U1884 ( .A0(n864), .A1(n2627), .B0(n185), .B1(n2629), .C0(n2626), 
        .Y(n1821) );
  AOI2BB2X1 U1885 ( .B0(stg2_real_7__7_), .B1(n875), .A0N(n858), .A1N(n2631), 
        .Y(n2626) );
  OAI221XL U1886 ( .A0(n864), .A1(n2636), .B0(n202), .B1(n2638), .C0(n2635), 
        .Y(n1822) );
  AOI2BB2X1 U1887 ( .B0(stg2_real_7__6_), .B1(n875), .A0N(n858), .A1N(n2640), 
        .Y(n2635) );
  OAI221XL U1888 ( .A0(n864), .A1(n2645), .B0(n203), .B1(n2647), .C0(n2644), 
        .Y(n1823) );
  AOI2BB2X1 U1889 ( .B0(stg2_real_7__5_), .B1(n869), .A0N(n857), .A1N(n2649), 
        .Y(n2644) );
  OAI221XL U1890 ( .A0(n864), .A1(n2654), .B0(n183), .B1(n2656), .C0(n2653), 
        .Y(n1824) );
  AOI2BB2X1 U1891 ( .B0(stg2_real_7__4_), .B1(n875), .A0N(n857), .A1N(n2658), 
        .Y(n2653) );
  OAI221XL U1892 ( .A0(n865), .A1(n2663), .B0(n195), .B1(n2665), .C0(n2662), 
        .Y(n1825) );
  AOI2BB2X1 U1893 ( .B0(stg2_real_7__3_), .B1(n869), .A0N(n857), .A1N(n2667), 
        .Y(n2662) );
  OAI221XL U1894 ( .A0(n865), .A1(n2672), .B0(n199), .B1(n2674), .C0(n2671), 
        .Y(n1826) );
  AOI2BB2X1 U1895 ( .B0(stg2_real_7__2_), .B1(n875), .A0N(n857), .A1N(n2676), 
        .Y(n2671) );
  OAI221XL U1896 ( .A0(n863), .A1(n2681), .B0(n185), .B1(n2683), .C0(n2680), 
        .Y(n1827) );
  AOI2BB2X1 U1897 ( .B0(stg2_real_7__1_), .B1(n875), .A0N(n857), .A1N(n2685), 
        .Y(n2680) );
  OAI221XL U1898 ( .A0(n9330), .A1(n2508), .B0(n853), .B1(n2970), .C0(n2506), 
        .Y(n1869) );
  AOI2BB2X1 U1899 ( .B0(stg2_img_15__7_), .B1(n872), .A0N(n2965), .A1N(n851), 
        .Y(n2506) );
  XOR2X1 U1900 ( .A(n3201), .B(n7430), .Y(stg2_img_15__7_) );
  OAI221XL U1901 ( .A0(n7270), .A1(n2514), .B0(n853), .B1(n2983), .C0(n2512), 
        .Y(n1870) );
  AOI2BB2X1 U1902 ( .B0(stg2_img_15__6_), .B1(n874), .A0N(n2978), .A1N(n852), 
        .Y(n2512) );
  XOR2X1 U1903 ( .A(n3200), .B(n7420), .Y(stg2_img_15__6_) );
  OAI221XL U1904 ( .A0(n9290), .A1(n2520), .B0(n853), .B1(n2996), .C0(n2518), 
        .Y(n1871) );
  XOR2X1 U1905 ( .A(n3199), .B(n7410), .Y(stg2_img_15__5_) );
  OAI221XL U1906 ( .A0(n7270), .A1(n2526), .B0(n854), .B1(n3009), .C0(n2524), 
        .Y(n1872) );
  XOR2X1 U1907 ( .A(n3198), .B(n7400), .Y(stg2_img_15__4_) );
  OAI221XL U1908 ( .A0(n9330), .A1(n2532), .B0(n853), .B1(n3022), .C0(n2530), 
        .Y(n1873) );
  AOI2BB2X1 U1909 ( .B0(stg2_img_15__3_), .B1(n873), .A0N(n3017), .A1N(n852), 
        .Y(n2530) );
  XOR2X1 U1910 ( .A(n3197), .B(n7390), .Y(stg2_img_15__3_) );
  OAI221XL U1911 ( .A0(n9330), .A1(n2538), .B0(n853), .B1(n3035), .C0(n2536), 
        .Y(n1874) );
  AOI2BB2X1 U1912 ( .B0(stg2_img_15__2_), .B1(n873), .A0N(n3030), .A1N(n852), 
        .Y(n2536) );
  XOR2X1 U1913 ( .A(n3196), .B(n7380), .Y(stg2_img_15__2_) );
  OAI221XL U1914 ( .A0(n9330), .A1(n2544), .B0(n853), .B1(n3048), .C0(n2542), 
        .Y(n1875) );
  AOI2BB2X1 U1915 ( .B0(stg2_img_15__1_), .B1(n873), .A0N(n3043), .A1N(n852), 
        .Y(n2542) );
  XOR2X1 U1916 ( .A(n3195), .B(n3194), .Y(stg2_img_15__1_) );
  OAI221XL U1917 ( .A0(n9330), .A1(n2638), .B0(n853), .B1(n2795), .C0(n2633), 
        .Y(n1854) );
  OAI221XL U1918 ( .A0(n9340), .A1(n2647), .B0(n853), .B1(n2805), .C0(n2642), 
        .Y(n1855) );
  OAI221XL U1919 ( .A0(n9340), .A1(n2656), .B0(n853), .B1(n2815), .C0(n2651), 
        .Y(n1856) );
  OAI221XL U1920 ( .A0(n9340), .A1(n2665), .B0(n853), .B1(n2825), .C0(n2660), 
        .Y(n1857) );
  AOI2BB1X1 U1921 ( .A0N(n2687), .A1N(n2663), .B0(n830), .Y(n2660) );
  OAI221XL U1922 ( .A0(n9340), .A1(n2674), .B0(n853), .B1(n2835), .C0(n2669), 
        .Y(n1858) );
  AOI2BB1X1 U1923 ( .A0N(n851), .A1N(n2672), .B0(n835), .Y(n2669) );
  OAI221XL U1924 ( .A0(n9340), .A1(n2683), .B0(n853), .B1(n2845), .C0(n2678), 
        .Y(n1859) );
  AOI2BB1X1 U1925 ( .A0N(n851), .A1N(n2681), .B0(n836), .Y(n2678) );
  OAI221XL U1926 ( .A0(n9340), .A1(n2694), .B0(n853), .B1(n2855), .C0(n2688), 
        .Y(n1860) );
  AOI2BB1X1 U1927 ( .A0N(n2692), .A1N(n852), .B0(n166), .Y(n2688) );
  OAI221XL U1928 ( .A0(n9330), .A1(n2550), .B0(n853), .B1(n3062), .C0(n2548), 
        .Y(n2308) );
  AOI2BB1X1 U1929 ( .A0N(n3057), .A1N(n852), .B0(n792), .Y(n2548) );
  OAI221XL U1930 ( .A0(n200), .A1(n2335), .B0(n82), .B1(n2627), .C0(n2333), 
        .Y(n2012) );
  AOI2BB2X1 U1931 ( .B0(stg2_real_5__7_), .B1(n872), .A0N(n850), .A1N(n2786), 
        .Y(n2333) );
  OAI221XL U1932 ( .A0(n189), .A1(n2342), .B0(n77), .B1(n2636), .C0(n2340), 
        .Y(n2013) );
  AOI2BB2X1 U1933 ( .B0(stg2_real_5__6_), .B1(n870), .A0N(n850), .A1N(n2796), 
        .Y(n2340) );
  OAI221XL U1934 ( .A0(n207), .A1(n2349), .B0(n80), .B1(n2645), .C0(n2347), 
        .Y(n2014) );
  AOI2BB2X1 U1935 ( .B0(stg2_real_5__5_), .B1(n870), .A0N(n850), .A1N(n2806), 
        .Y(n2347) );
  OAI221XL U1936 ( .A0(n197), .A1(n2356), .B0(n76), .B1(n2654), .C0(n2354), 
        .Y(n2015) );
  AOI2BB2X1 U1937 ( .B0(stg2_real_5__4_), .B1(n870), .A0N(n850), .A1N(n2816), 
        .Y(n2354) );
  OAI221XL U1938 ( .A0(n200), .A1(n2363), .B0(n75), .B1(n2663), .C0(n2361), 
        .Y(n2016) );
  AOI2BB2X1 U1939 ( .B0(stg2_real_5__3_), .B1(n870), .A0N(n850), .A1N(n2826), 
        .Y(n2361) );
  OAI221XL U1940 ( .A0(n202), .A1(n2370), .B0(n75), .B1(n2672), .C0(n2368), 
        .Y(n2017) );
  AOI2BB2X1 U1941 ( .B0(stg2_real_5__2_), .B1(n871), .A0N(n850), .A1N(n2836), 
        .Y(n2368) );
  OAI221XL U1942 ( .A0(n203), .A1(n2377), .B0(n76), .B1(n2681), .C0(n2375), 
        .Y(n2018) );
  AOI2BB2X1 U1943 ( .B0(stg2_real_5__1_), .B1(n874), .A0N(n850), .A1N(n2846), 
        .Y(n2375) );
  OAI221XL U1944 ( .A0(n205), .A1(n2384), .B0(n79), .B1(n2692), .C0(n2382), 
        .Y(n2019) );
  AOI2BB2X1 U1945 ( .B0(stg2_real_5__0_), .B1(n871), .A0N(n850), .A1N(n2856), 
        .Y(n2382) );
  OAI221XL U1946 ( .A0(n906), .A1(n2692), .B0(n46), .B1(n1413), .C0(n1410), 
        .Y(n1987) );
  AOI2BB1X1 U1947 ( .A0N(n902), .A1N(n98), .B0(n165), .Y(n1410) );
  OAI221XL U1948 ( .A0(n917), .A1(n2692), .B0(n50), .B1(n2694), .C0(n2689), 
        .Y(n1891) );
  AOI2BB1X1 U1949 ( .A0N(n856), .A1N(n2851), .B0(n166), .Y(n2689) );
  OAI221XL U1950 ( .A0(n908), .A1(n2618), .B0(n49), .B1(n1349), .C0(n1346), 
        .Y(n1979) );
  AOI2BB1X1 U1951 ( .A0N(n902), .A1N(n124), .B0(n814), .Y(n1346) );
  OAI221XL U1952 ( .A0(n908), .A1(n2627), .B0(n45), .B1(n1357), .C0(n1354), 
        .Y(n1980) );
  AOI2BB1X1 U1953 ( .A0N(n902), .A1N(n125), .B0(n815), .Y(n1354) );
  OAI221XL U1954 ( .A0(n908), .A1(n2636), .B0(n52), .B1(n1365), .C0(n1362), 
        .Y(n1981) );
  AOI2BB1X1 U1955 ( .A0N(n902), .A1N(n126), .B0(n816), .Y(n1362) );
  OAI221XL U1956 ( .A0(n906), .A1(n2645), .B0(n19), .B1(n1373), .C0(n1370), 
        .Y(n1982) );
  AOI2BB1X1 U1957 ( .A0N(n902), .A1N(n117), .B0(n817), .Y(n1370) );
  OAI221XL U1958 ( .A0(n906), .A1(n2654), .B0(n20), .B1(n1381), .C0(n1378), 
        .Y(n1983) );
  AOI2BB1X1 U1959 ( .A0N(n902), .A1N(n118), .B0(n818), .Y(n1378) );
  OAI221XL U1960 ( .A0(n907), .A1(n2663), .B0(n49), .B1(n1389), .C0(n1386), 
        .Y(n1984) );
  AOI2BB1X1 U1961 ( .A0N(n902), .A1N(n119), .B0(n819), .Y(n1386) );
  OAI221XL U1962 ( .A0(n907), .A1(n2672), .B0(n45), .B1(n1397), .C0(n1394), 
        .Y(n1985) );
  AOI2BB1X1 U1963 ( .A0N(n902), .A1N(n115), .B0(n820), .Y(n1394) );
  OAI221XL U1964 ( .A0(n906), .A1(n2681), .B0(n46), .B1(n1405), .C0(n1402), 
        .Y(n1986) );
  AOI2BB1X1 U1965 ( .A0N(n902), .A1N(n116), .B0(n821), .Y(n1402) );
  OAI221XL U1966 ( .A0(n917), .A1(n2618), .B0(n49), .B1(n2620), .C0(n2616), 
        .Y(n1883) );
  AOI2BB1X1 U1967 ( .A0N(n856), .A1N(n2771), .B0(n825), .Y(n2616) );
  OAI221XL U1968 ( .A0(n9200), .A1(n2627), .B0(n52), .B1(n2629), .C0(n2625), 
        .Y(n1884) );
  AOI2BB1X1 U1969 ( .A0N(n856), .A1N(n2781), .B0(n826), .Y(n2625) );
  OAI221XL U1970 ( .A0(n917), .A1(n2636), .B0(n45), .B1(n2638), .C0(n2634), 
        .Y(n1885) );
  AOI2BB1X1 U1971 ( .A0N(n856), .A1N(n2791), .B0(n827), .Y(n2634) );
  OAI221XL U1972 ( .A0(n917), .A1(n2645), .B0(n47), .B1(n2647), .C0(n2643), 
        .Y(n1886) );
  AOI2BB1X1 U1973 ( .A0N(n856), .A1N(n2801), .B0(n828), .Y(n2643) );
  OAI221XL U1974 ( .A0(n917), .A1(n2654), .B0(n46), .B1(n2656), .C0(n2652), 
        .Y(n1887) );
  AOI2BB1X1 U1975 ( .A0N(n856), .A1N(n2811), .B0(n829), .Y(n2652) );
  OAI221XL U1976 ( .A0(n917), .A1(n2663), .B0(n48), .B1(n2665), .C0(n2661), 
        .Y(n1888) );
  AOI2BB1X1 U1977 ( .A0N(n856), .A1N(n2821), .B0(n830), .Y(n2661) );
  OAI221XL U1978 ( .A0(n917), .A1(n2672), .B0(n48), .B1(n2674), .C0(n2670), 
        .Y(n1889) );
  AOI2BB1X1 U1979 ( .A0N(n856), .A1N(n2831), .B0(n835), .Y(n2670) );
  OAI221XL U1980 ( .A0(n9190), .A1(n2681), .B0(n45), .B1(n2683), .C0(n2679), 
        .Y(n1890) );
  AOI2BB1X1 U1981 ( .A0N(n856), .A1N(n2841), .B0(n836), .Y(n2679) );
  OAI221XL U1982 ( .A0(n917), .A1(n3057), .B0(n49), .B1(n2550), .C0(n2549), 
        .Y(n1907) );
  AOI2BB1X1 U1983 ( .A0N(n856), .A1N(n3059), .B0(n792), .Y(n2549) );
  OAI221XL U1984 ( .A0(n909), .A1(n3057), .B0(n45), .B1(n3058), .C0(n3054), 
        .Y(n2003) );
  AOI2BB1X1 U1985 ( .A0N(n902), .A1N(n114), .B0(n793), .Y(n3054) );
  OAI221XL U1986 ( .A0(n2953), .A1(n9310), .B0(n9270), .B1(n2952), .C0(n2951), 
        .Y(n1963) );
  AOI2BB2X1 U1987 ( .B0(stg2_img_14__8_), .B1(n869), .A0N(n9230), .A1N(n3111), 
        .Y(n2951) );
  XOR2X1 U1988 ( .A(n3189), .B(n7680), .Y(stg2_img_14__8_) );
  OAI221XL U1989 ( .A0(n2966), .A1(n9350), .B0(n9270), .B1(n2965), .C0(n2964), 
        .Y(n1964) );
  AOI2BB2X1 U1990 ( .B0(stg2_img_14__7_), .B1(n875), .A0N(n9230), .A1N(n3115), 
        .Y(n2964) );
  XOR2X1 U1991 ( .A(n3188), .B(n7530), .Y(stg2_img_14__7_) );
  OAI221XL U1992 ( .A0(n2979), .A1(n9320), .B0(n9270), .B1(n2978), .C0(n2977), 
        .Y(n1965) );
  AOI2BB2X1 U1993 ( .B0(stg2_img_14__6_), .B1(n870), .A0N(n9230), .A1N(n3120), 
        .Y(n2977) );
  XOR2X1 U1994 ( .A(n3187), .B(n7650), .Y(stg2_img_14__6_) );
  OAI221XL U1995 ( .A0(n2992), .A1(n9310), .B0(n9270), .B1(n2991), .C0(n2990), 
        .Y(n1966) );
  AOI2BB2X1 U1996 ( .B0(stg2_img_14__5_), .B1(n869), .A0N(n9230), .A1N(n3125), 
        .Y(n2990) );
  XOR2X1 U1997 ( .A(n3186), .B(n7500), .Y(stg2_img_14__5_) );
  OAI221XL U1998 ( .A0(n3005), .A1(n9290), .B0(n9270), .B1(n3004), .C0(n3003), 
        .Y(n1967) );
  AOI2BB2X1 U1999 ( .B0(stg2_img_14__4_), .B1(n870), .A0N(n9230), .A1N(n3129), 
        .Y(n3003) );
  XOR2X1 U2000 ( .A(n3185), .B(n7620), .Y(stg2_img_14__4_) );
  OAI221XL U2001 ( .A0(n3018), .A1(n9300), .B0(n9270), .B1(n3017), .C0(n3016), 
        .Y(n1968) );
  AOI2BB2X1 U2002 ( .B0(stg2_img_14__3_), .B1(n869), .A0N(n9230), .A1N(n3133), 
        .Y(n3016) );
  XOR2X1 U2003 ( .A(n3184), .B(n7590), .Y(stg2_img_14__3_) );
  OAI221XL U2004 ( .A0(n3031), .A1(n9320), .B0(n9270), .B1(n3030), .C0(n3029), 
        .Y(n1969) );
  AOI2BB2X1 U2005 ( .B0(stg2_img_14__2_), .B1(n869), .A0N(n9230), .A1N(n3137), 
        .Y(n3029) );
  XOR2X1 U2006 ( .A(n3183), .B(n7560), .Y(stg2_img_14__2_) );
  OAI221XL U2007 ( .A0(n3044), .A1(n9300), .B0(n9260), .B1(n3043), .C0(n3042), 
        .Y(n1970) );
  AOI2BB2X1 U2008 ( .B0(stg2_img_14__1_), .B1(n869), .A0N(n9230), .A1N(n3141), 
        .Y(n3042) );
  XOR2X1 U2009 ( .A(n3182), .B(n3181), .Y(stg2_img_14__1_) );
  OAI221XL U2010 ( .A0(n3058), .A1(n9320), .B0(n9270), .B1(n3057), .C0(n3056), 
        .Y(n1971) );
  AOI2BB1X1 U2011 ( .A0N(n9240), .A1N(n3147), .B0(n793), .Y(n3056) );
  OAI221XL U2012 ( .A0(n50), .A1(n2328), .B0(n207), .B1(n2618), .C0(n2325), 
        .Y(n2075) );
  AOI2BB1X1 U2013 ( .A0N(n848), .A1N(n2773), .B0(n800), .Y(n2325) );
  OAI221XL U2014 ( .A0(n9290), .A1(n1349), .B0(n9260), .B1(n2618), .C0(n1345), 
        .Y(n1947) );
  AOI2BB1X1 U2015 ( .A0N(n3079), .A1N(n2772), .B0(n814), .Y(n1345) );
  OAI221XL U2016 ( .A0(n9310), .A1(n1357), .B0(n9260), .B1(n2627), .C0(n1353), 
        .Y(n1948) );
  AOI2BB1X1 U2017 ( .A0N(n3079), .A1N(n2782), .B0(n815), .Y(n1353) );
  OAI221XL U2018 ( .A0(n9300), .A1(n1365), .B0(n9260), .B1(n2636), .C0(n1361), 
        .Y(n1949) );
  AOI2BB1X1 U2019 ( .A0N(n9240), .A1N(n2792), .B0(n816), .Y(n1361) );
  OAI221XL U2020 ( .A0(n9320), .A1(n1373), .B0(n9260), .B1(n2645), .C0(n1369), 
        .Y(n1950) );
  AOI2BB1X1 U2021 ( .A0N(n9240), .A1N(n2802), .B0(n817), .Y(n1369) );
  OAI221XL U2022 ( .A0(n9310), .A1(n1381), .B0(n9260), .B1(n2654), .C0(n1377), 
        .Y(n1951) );
  AOI2BB1X1 U2023 ( .A0N(n9240), .A1N(n2812), .B0(n818), .Y(n1377) );
  OAI221XL U2024 ( .A0(n9310), .A1(n1389), .B0(n9260), .B1(n2663), .C0(n1385), 
        .Y(n1952) );
  AOI2BB1X1 U2025 ( .A0N(n9240), .A1N(n2822), .B0(n819), .Y(n1385) );
  OAI221XL U2026 ( .A0(n9350), .A1(n1397), .B0(n9260), .B1(n2672), .C0(n1393), 
        .Y(n1953) );
  AOI2BB1X1 U2027 ( .A0N(n9240), .A1N(n2832), .B0(n820), .Y(n1393) );
  OAI221XL U2028 ( .A0(n9330), .A1(n1405), .B0(n9270), .B1(n2681), .C0(n1401), 
        .Y(n1954) );
  AOI2BB1X1 U2029 ( .A0N(n9240), .A1N(n2842), .B0(n821), .Y(n1401) );
  OAI221XL U2030 ( .A0(n9320), .A1(n1413), .B0(n9270), .B1(n2692), .C0(n1409), 
        .Y(n1955) );
  AOI2BB1X1 U2031 ( .A0N(n9240), .A1N(n2852), .B0(n165), .Y(n1409) );
  OAI221XL U2032 ( .A0(n9310), .A1(n2328), .B0(n45), .B1(n2618), .C0(n2324), 
        .Y(n2043) );
  AOI2BB1X1 U2033 ( .A0N(n2456), .A1N(n2774), .B0(n800), .Y(n2324) );
  OAI221XL U2034 ( .A0(n49), .A1(n2335), .B0(n185), .B1(n2627), .C0(n2332), 
        .Y(n2076) );
  AOI2BB1X1 U2035 ( .A0N(n848), .A1N(n2783), .B0(n801), .Y(n2332) );
  OAI221XL U2036 ( .A0(n9310), .A1(n2335), .B0(n50), .B1(n2627), .C0(n2331), 
        .Y(n2044) );
  AOI2BB1X1 U2037 ( .A0N(n846), .A1N(n2784), .B0(n801), .Y(n2331) );
  OAI221XL U2038 ( .A0(n19), .A1(n2342), .B0(n189), .B1(n2636), .C0(n2339), 
        .Y(n2077) );
  AOI2BB1X1 U2039 ( .A0N(n848), .A1N(n2793), .B0(n802), .Y(n2339) );
  OAI221XL U2040 ( .A0(n9310), .A1(n2342), .B0(n20), .B1(n2636), .C0(n2338), 
        .Y(n2045) );
  AOI2BB1X1 U2041 ( .A0N(n846), .A1N(n2794), .B0(n802), .Y(n2338) );
  OAI221XL U2042 ( .A0(n20), .A1(n2349), .B0(n197), .B1(n2645), .C0(n2346), 
        .Y(n2078) );
  AOI2BB1X1 U2043 ( .A0N(n848), .A1N(n2803), .B0(n803), .Y(n2346) );
  OAI221XL U2044 ( .A0(n9310), .A1(n2349), .B0(n20), .B1(n2645), .C0(n2345), 
        .Y(n2046) );
  AOI2BB1X1 U2045 ( .A0N(n846), .A1N(n2804), .B0(n803), .Y(n2345) );
  OAI221XL U2046 ( .A0(n46), .A1(n2356), .B0(n187), .B1(n2654), .C0(n2353), 
        .Y(n2079) );
  AOI2BB1X1 U2047 ( .A0N(n848), .A1N(n2813), .B0(n804), .Y(n2353) );
  OAI221XL U2048 ( .A0(n9310), .A1(n2356), .B0(n46), .B1(n2654), .C0(n2352), 
        .Y(n2047) );
  AOI2BB1X1 U2049 ( .A0N(n846), .A1N(n2814), .B0(n804), .Y(n2352) );
  OAI221XL U2050 ( .A0(n52), .A1(n2363), .B0(n200), .B1(n2663), .C0(n2360), 
        .Y(n2080) );
  AOI2BB1X1 U2051 ( .A0N(n848), .A1N(n2823), .B0(n805), .Y(n2360) );
  OAI221XL U2052 ( .A0(n9320), .A1(n2363), .B0(n47), .B1(n2663), .C0(n2359), 
        .Y(n2048) );
  AOI2BB1X1 U2053 ( .A0N(n846), .A1N(n2824), .B0(n805), .Y(n2359) );
  OAI221XL U2054 ( .A0(n45), .A1(n2370), .B0(n187), .B1(n2672), .C0(n2367), 
        .Y(n2081) );
  AOI2BB1X1 U2055 ( .A0N(n848), .A1N(n2833), .B0(n806), .Y(n2367) );
  OAI221XL U2056 ( .A0(n9310), .A1(n2370), .B0(n51), .B1(n2672), .C0(n2366), 
        .Y(n2049) );
  AOI2BB1X1 U2057 ( .A0N(n846), .A1N(n2834), .B0(n806), .Y(n2366) );
  OAI221XL U2058 ( .A0(n50), .A1(n2377), .B0(n207), .B1(n2681), .C0(n2374), 
        .Y(n2082) );
  AOI2BB1X1 U2059 ( .A0N(n848), .A1N(n2843), .B0(n807), .Y(n2374) );
  OAI221XL U2060 ( .A0(n9310), .A1(n2377), .B0(n49), .B1(n2681), .C0(n2373), 
        .Y(n2050) );
  AOI2BB1X1 U2061 ( .A0N(n846), .A1N(n2844), .B0(n807), .Y(n2373) );
  OAI221XL U2062 ( .A0(n51), .A1(n2384), .B0(n185), .B1(n2692), .C0(n2381), 
        .Y(n2083) );
  AOI2BB1X1 U2063 ( .A0N(n848), .A1N(n2853), .B0(n167), .Y(n2381) );
  OAI221XL U2064 ( .A0(n9310), .A1(n2384), .B0(n47), .B1(n2692), .C0(n2380), 
        .Y(n2051) );
  AOI2BB1X1 U2065 ( .A0N(n846), .A1N(n2854), .B0(n167), .Y(n2380) );
  OAI221XL U2066 ( .A0(n9320), .A1(n2418), .B0(n48), .B1(n2952), .C0(n2416), 
        .Y(n2059) );
  AOI2BB2X1 U2067 ( .B0(stg2_img_13__8_), .B1(n872), .A0N(n845), .A1N(n2956), 
        .Y(n2416) );
  XOR2X1 U2068 ( .A(n3174), .B(n7690), .Y(stg2_img_13__8_) );
  OAI221XL U2069 ( .A0(n9350), .A1(n2423), .B0(n19), .B1(n2965), .C0(n2421), 
        .Y(n2060) );
  AOI2BB2X1 U2070 ( .B0(stg2_img_13__7_), .B1(n871), .A0N(n845), .A1N(n2969), 
        .Y(n2421) );
  XOR2X1 U2071 ( .A(n3173), .B(n7540), .Y(stg2_img_13__7_) );
  OAI221XL U2072 ( .A0(n9320), .A1(n2428), .B0(n52), .B1(n2978), .C0(n2426), 
        .Y(n2061) );
  AOI2BB2X1 U2073 ( .B0(stg2_img_13__6_), .B1(n871), .A0N(n845), .A1N(n2982), 
        .Y(n2426) );
  XOR2X1 U2074 ( .A(n3172), .B(n7660), .Y(stg2_img_13__6_) );
  OAI221XL U2075 ( .A0(n9290), .A1(n2433), .B0(n51), .B1(n2991), .C0(n2431), 
        .Y(n2062) );
  AOI2BB2X1 U2076 ( .B0(stg2_img_13__5_), .B1(n871), .A0N(n845), .A1N(n2995), 
        .Y(n2431) );
  XOR2X1 U2077 ( .A(n3171), .B(n7510), .Y(stg2_img_13__5_) );
  OAI221XL U2078 ( .A0(n9320), .A1(n2438), .B0(n19), .B1(n3004), .C0(n2436), 
        .Y(n2063) );
  AOI2BB2X1 U2079 ( .B0(stg2_img_13__4_), .B1(n871), .A0N(n845), .A1N(n3008), 
        .Y(n2436) );
  XOR2X1 U2080 ( .A(n3170), .B(n7630), .Y(stg2_img_13__4_) );
  OAI221XL U2081 ( .A0(n9290), .A1(n2443), .B0(n46), .B1(n3017), .C0(n2441), 
        .Y(n2064) );
  AOI2BB2X1 U2082 ( .B0(stg2_img_13__3_), .B1(n871), .A0N(n845), .A1N(n3021), 
        .Y(n2441) );
  XOR2X1 U2083 ( .A(n3169), .B(n7600), .Y(stg2_img_13__3_) );
  OAI221XL U2084 ( .A0(n9320), .A1(n2448), .B0(n51), .B1(n3030), .C0(n2446), 
        .Y(n2065) );
  AOI2BB2X1 U2085 ( .B0(stg2_img_13__2_), .B1(n871), .A0N(n845), .A1N(n3034), 
        .Y(n2446) );
  XOR2X1 U2086 ( .A(n3168), .B(n7570), .Y(stg2_img_13__2_) );
  OAI221XL U2087 ( .A0(n9320), .A1(n2453), .B0(n52), .B1(n3043), .C0(n2451), 
        .Y(n2066) );
  AOI2BB2X1 U2088 ( .B0(stg2_img_13__1_), .B1(n871), .A0N(n845), .A1N(n3047), 
        .Y(n2451) );
  XOR2X1 U2089 ( .A(n3167), .B(n3166), .Y(stg2_img_13__1_) );
  OAI221XL U2090 ( .A0(n52), .A1(n2461), .B0(n181), .B1(n3057), .C0(n2459), 
        .Y(n2099) );
  AOI2BB1X1 U2091 ( .A0N(n848), .A1N(n3060), .B0(n831), .Y(n2459) );
  OAI221XL U2092 ( .A0(n9320), .A1(n2461), .B0(n19), .B1(n3057), .C0(n2457), 
        .Y(n2067) );
  AOI2BB1X1 U2093 ( .A0N(n846), .A1N(n3061), .B0(n831), .Y(n2457) );
  OAI221XL U2094 ( .A0(n855), .A1(n2967), .B0(n892), .B1(n3201), .C0(n2507), 
        .Y(n1900) );
  OAI221XL U2095 ( .A0(n855), .A1(n2980), .B0(n891), .B1(n3200), .C0(n2513), 
        .Y(n1901) );
  OAI221XL U2096 ( .A0(n855), .A1(n2993), .B0(n891), .B1(n3199), .C0(n2519), 
        .Y(n1902) );
  OAI221XL U2097 ( .A0(n855), .A1(n3006), .B0(n891), .B1(n3198), .C0(n2525), 
        .Y(n1903) );
  OAI221XL U2098 ( .A0(n856), .A1(n3019), .B0(n891), .B1(n3197), .C0(n2531), 
        .Y(n1904) );
  OAI221XL U2099 ( .A0(n856), .A1(n3032), .B0(n891), .B1(n3196), .C0(n2537), 
        .Y(n1905) );
  OAI221XL U2100 ( .A0(n856), .A1(n3045), .B0(n890), .B1(n3195), .C0(n2543), 
        .Y(n1906) );
  OAI221XL U2101 ( .A0(n901), .A1(n101), .B0(n890), .B1(n3185), .C0(n3002), 
        .Y(n1999) );
  OA22X1 U2102 ( .A0(n908), .A1(n3004), .B0(n19), .B1(n3005), .Y(n3002) );
  OAI221XL U2103 ( .A0(n901), .A1(n99), .B0(n888), .B1(n3183), .C0(n3028), .Y(
        n2001) );
  OA22X1 U2104 ( .A0(n908), .A1(n3030), .B0(n45), .B1(n3031), .Y(n3028) );
  OAI221XL U2105 ( .A0(n901), .A1(n100), .B0(n893), .B1(n3182), .C0(n3041), 
        .Y(n2002) );
  OA22X1 U2106 ( .A0(n908), .A1(n3043), .B0(n51), .B1(n3044), .Y(n3041) );
  OAI221XL U2107 ( .A0(n847), .A1(n2968), .B0(n894), .B1(n3173), .C0(n2422), 
        .Y(n2092) );
  OAI221XL U2108 ( .A0(n847), .A1(n2981), .B0(n894), .B1(n3172), .C0(n2427), 
        .Y(n2093) );
  OAI221XL U2109 ( .A0(n847), .A1(n2994), .B0(n894), .B1(n3171), .C0(n2432), 
        .Y(n2094) );
  OAI221XL U2110 ( .A0(n847), .A1(n3007), .B0(n894), .B1(n3170), .C0(n2437), 
        .Y(n2095) );
  OAI221XL U2111 ( .A0(n847), .A1(n3020), .B0(n894), .B1(n3169), .C0(n2442), 
        .Y(n2096) );
  OAI221XL U2112 ( .A0(n847), .A1(n3033), .B0(n893), .B1(n3168), .C0(n2447), 
        .Y(n2097) );
  OAI221XL U2113 ( .A0(n847), .A1(n3046), .B0(n893), .B1(n3167), .C0(n2452), 
        .Y(n2098) );
  OAI221XL U2114 ( .A0(n901), .A1(n105), .B0(n889), .B1(n3188), .C0(n2963), 
        .Y(n1996) );
  OAI221XL U2115 ( .A0(n901), .A1(n3119), .B0(n889), .B1(n3187), .C0(n2976), 
        .Y(n1997) );
  OAI221XL U2116 ( .A0(n901), .A1(n3124), .B0(n889), .B1(n3186), .C0(n2989), 
        .Y(n1998) );
  OA22X1 U2117 ( .A0(n908), .A1(n2991), .B0(n50), .B1(n2992), .Y(n2989) );
  OAI221XL U2118 ( .A0(n901), .A1(n102), .B0(n888), .B1(n3184), .C0(n3015), 
        .Y(n2000) );
  OA22X1 U2119 ( .A0(n908), .A1(n3017), .B0(n52), .B1(n3018), .Y(n3015) );
  OA22X1 U2120 ( .A0(n199), .A1(n1280), .B0(n82), .B1(n1279), .Y(n1281) );
  OA22X1 U2121 ( .A0(n185), .A1(n2685), .B0(n77), .B1(n2684), .Y(n2686) );
  OA22X1 U2122 ( .A0(n183), .A1(n2676), .B0(n78), .B1(n2675), .Y(n2677) );
  OA22X1 U2123 ( .A0(n181), .A1(n2667), .B0(n84), .B1(n2666), .Y(n2668) );
  OA22X1 U2124 ( .A0(n195), .A1(n2658), .B0(n83), .B1(n2657), .Y(n2659) );
  OA22X1 U2125 ( .A0(n205), .A1(n2649), .B0(n84), .B1(n2648), .Y(n2650) );
  OA22X1 U2126 ( .A0(n207), .A1(n2640), .B0(n80), .B1(n2639), .Y(n2641) );
  OA22X1 U2127 ( .A0(n187), .A1(n2631), .B0(n76), .B1(n2630), .Y(n2632) );
  OA22X1 U2128 ( .A0(n187), .A1(n2622), .B0(n76), .B1(n2621), .Y(n2623) );
  OA22X1 U2129 ( .A0(n203), .A1(n1407), .B0(n81), .B1(n1406), .Y(n1408) );
  OA22X1 U2130 ( .A0(n200), .A1(n1399), .B0(n80), .B1(n1398), .Y(n1400) );
  OA22X1 U2131 ( .A0(n202), .A1(n1391), .B0(n77), .B1(n1390), .Y(n1392) );
  OA22X1 U2132 ( .A0(n181), .A1(n1383), .B0(n75), .B1(n1382), .Y(n1384) );
  OA22X1 U2133 ( .A0(n195), .A1(n1375), .B0(n83), .B1(n1374), .Y(n1376) );
  OA22X1 U2134 ( .A0(n203), .A1(n1367), .B0(n81), .B1(n1366), .Y(n1368) );
  OA22X1 U2135 ( .A0(n195), .A1(n1359), .B0(n80), .B1(n1358), .Y(n1360) );
  OAI221X1 U2136 ( .A0(n9760), .A1(n2852), .B0(n48), .B1(n98), .C0(n1416), .Y(
        stg2_real_Wn[16]) );
  OA22X1 U2137 ( .A0(n205), .A1(n1415), .B0(n79), .B1(n1414), .Y(n1416) );
  OA22X1 U2138 ( .A0(n203), .A1(n1271), .B0(n77), .B1(n1270), .Y(n1272) );
  OA22X1 U2139 ( .A0(n195), .A1(n1262), .B0(n76), .B1(n1261), .Y(n1263) );
  OA22X1 U2140 ( .A0(n200), .A1(n1253), .B0(n82), .B1(n1252), .Y(n1254) );
  OA22X1 U2141 ( .A0(n203), .A1(n1244), .B0(n79), .B1(n1243), .Y(n1245) );
  OA22X1 U2142 ( .A0(n197), .A1(n1235), .B0(n76), .B1(n1234), .Y(n1236) );
  OA22X1 U2143 ( .A0(n199), .A1(n1226), .B0(n75), .B1(n1225), .Y(n1227) );
  OA22X1 U2144 ( .A0(n199), .A1(n2846), .B0(n84), .B1(n2378), .Y(n2379) );
  OA22X1 U2145 ( .A0(n181), .A1(n2836), .B0(n84), .B1(n2371), .Y(n2372) );
  OA22X1 U2146 ( .A0(n189), .A1(n2826), .B0(n83), .B1(n2364), .Y(n2365) );
  OAI222XL U2147 ( .A0(n898), .A1(n3165), .B0(n7330), .B1(n10620), .C0(n52), 
        .C1(n10550), .Y(n2164) );
  OAI222XL U2148 ( .A0(n123), .A1(n891), .B0(n7340), .B1(n10630), .C0(n9300), 
        .C1(n10550), .Y(n2132) );
  CLKINVX1 U2149 ( .A(stg2_img_8__15_), .Y(n3165) );
  OAI222XL U2150 ( .A0(n898), .A1(n3164), .B0(n7330), .B1(n10670), .C0(n47), 
        .C1(n10640), .Y(n2165) );
  OAI222XL U2151 ( .A0(n121), .A1(n898), .B0(n7340), .B1(n10680), .C0(n9300), 
        .C1(n10640), .Y(n2133) );
  OAI222XL U2152 ( .A0(n898), .A1(n3163), .B0(n7330), .B1(n10720), .C0(n49), 
        .C1(n10690), .Y(n2166) );
  OAI222XL U2153 ( .A0(n122), .A1(n897), .B0(n7340), .B1(n10730), .C0(n9300), 
        .C1(n10690), .Y(n2134) );
  OAI222XL U2154 ( .A0(n898), .A1(n3162), .B0(n7330), .B1(n10770), .C0(n48), 
        .C1(n10740), .Y(n2167) );
  OAI222XL U2155 ( .A0(n129), .A1(n891), .B0(n7340), .B1(n10780), .C0(n9300), 
        .C1(n10740), .Y(n2135) );
  OAI222XL U2156 ( .A0(n898), .A1(n3161), .B0(n7330), .B1(n10820), .C0(n45), 
        .C1(n10790), .Y(n2168) );
  OAI222XL U2157 ( .A0(n130), .A1(n898), .B0(n7340), .B1(n10830), .C0(n9300), 
        .C1(n10790), .Y(n2136) );
  OAI222XL U2158 ( .A0(n897), .A1(n3160), .B0(n7330), .B1(n10870), .C0(n46), 
        .C1(n10840), .Y(n2169) );
  OAI222XL U2159 ( .A0(n131), .A1(n896), .B0(n7340), .B1(n10880), .C0(n9300), 
        .C1(n10840), .Y(n2137) );
  OAI222XL U2160 ( .A0(n897), .A1(n3159), .B0(n7330), .B1(n10920), .C0(n48), 
        .C1(n10890), .Y(n2170) );
  OAI222XL U2161 ( .A0(n147), .A1(n895), .B0(n7340), .B1(n10930), .C0(n9300), 
        .C1(n10890), .Y(n2138) );
  OAI221XL U2162 ( .A0(n844), .A1(n2704), .B0(n205), .B1(n2702), .C0(n2699), 
        .Y(n3209) );
  NAND2X1 U2163 ( .A(stg2_real_4__15_), .B(n886), .Y(n2699) );
  OAI221XL U2164 ( .A0(n844), .A1(n1154), .B0(n207), .B1(n1152), .C0(n1150), 
        .Y(n3210) );
  NAND2X1 U2165 ( .A(stg2_real_4__14_), .B(n879), .Y(n1150) );
  OAI221XL U2166 ( .A0(n844), .A1(n1163), .B0(n183), .B1(n1161), .C0(n1159), 
        .Y(n3211) );
  NAND2X1 U2167 ( .A(stg2_real_4__13_), .B(n877), .Y(n1159) );
  OAI221XL U2168 ( .A0(n844), .A1(n1172), .B0(n205), .B1(n1170), .C0(n1168), 
        .Y(n3212) );
  NAND2X1 U2169 ( .A(stg2_real_4__12_), .B(n877), .Y(n1168) );
  OAI221XL U2170 ( .A0(n844), .A1(n1181), .B0(n200), .B1(n1179), .C0(n1177), 
        .Y(n3213) );
  NAND2X1 U2171 ( .A(stg2_real_4__11_), .B(n878), .Y(n1177) );
  OAI221XL U2172 ( .A0(n844), .A1(n1190), .B0(n197), .B1(n1188), .C0(n1186), 
        .Y(n3214) );
  NAND2X1 U2173 ( .A(stg2_real_4__10_), .B(n876), .Y(n1186) );
  OAI221XL U2174 ( .A0(n844), .A1(n1199), .B0(n187), .B1(n1197), .C0(n1195), 
        .Y(n3215) );
  NAND2X1 U2175 ( .A(stg2_real_4__9_), .B(n876), .Y(n1195) );
  OAI221XL U2176 ( .A0(n844), .A1(n1208), .B0(n185), .B1(n1206), .C0(n1204), 
        .Y(n3216) );
  NAND2X1 U2177 ( .A(stg2_real_4__8_), .B(n876), .Y(n1204) );
  OAI221XL U2178 ( .A0(n9380), .A1(n2703), .B0(n84), .B1(n2702), .C0(n2701), 
        .Y(n2180) );
  NAND2X1 U2179 ( .A(stg2_real_0__15_), .B(n878), .Y(n2701) );
  OAI221XL U2180 ( .A0(n7330), .A1(n2706), .B0(n51), .B1(n2702), .C0(n2698), 
        .Y(n2148) );
  OAI221XL U2181 ( .A0(n7340), .A1(n2707), .B0(n9330), .B1(n2702), .C0(n2698), 
        .Y(n2116) );
  OAI221XL U2182 ( .A0(n9360), .A1(n1153), .B0(n77), .B1(n1152), .C0(n1151), 
        .Y(n2181) );
  NAND2X1 U2183 ( .A(stg2_real_0__14_), .B(n877), .Y(n1151) );
  OAI221XL U2184 ( .A0(n860), .A1(n1156), .B0(n47), .B1(n1152), .C0(n1148), 
        .Y(n2149) );
  OAI221XL U2185 ( .A0(n859), .A1(n1157), .B0(n9290), .B1(n1152), .C0(n1148), 
        .Y(n2117) );
  OAI221XL U2186 ( .A0(n9360), .A1(n1162), .B0(n82), .B1(n1161), .C0(n1160), 
        .Y(n2182) );
  NAND2X1 U2187 ( .A(stg2_real_0__13_), .B(n877), .Y(n1160) );
  OAI221XL U2188 ( .A0(n860), .A1(n1165), .B0(n19), .B1(n1161), .C0(n1158), 
        .Y(n2150) );
  OAI221XL U2189 ( .A0(n859), .A1(n1166), .B0(n9290), .B1(n1161), .C0(n1158), 
        .Y(n2118) );
  OAI221XL U2190 ( .A0(n9360), .A1(n1171), .B0(n75), .B1(n1170), .C0(n1169), 
        .Y(n2183) );
  NAND2X1 U2191 ( .A(stg2_real_0__12_), .B(n877), .Y(n1169) );
  OAI221XL U2192 ( .A0(n860), .A1(n1174), .B0(n48), .B1(n1170), .C0(n1167), 
        .Y(n2151) );
  OAI221XL U2193 ( .A0(n859), .A1(n1175), .B0(n9340), .B1(n1170), .C0(n1167), 
        .Y(n2119) );
  OAI221XL U2194 ( .A0(n9360), .A1(n1180), .B0(n75), .B1(n1179), .C0(n1178), 
        .Y(n2184) );
  NAND2X1 U2195 ( .A(stg2_real_0__11_), .B(n878), .Y(n1178) );
  OAI221XL U2196 ( .A0(n860), .A1(n1183), .B0(n50), .B1(n1179), .C0(n1176), 
        .Y(n2152) );
  OAI221XL U2197 ( .A0(n859), .A1(n1184), .B0(n9290), .B1(n1179), .C0(n1176), 
        .Y(n2120) );
  OAI221XL U2198 ( .A0(n9360), .A1(n1189), .B0(n82), .B1(n1188), .C0(n1187), 
        .Y(n2185) );
  NAND2X1 U2199 ( .A(stg2_real_0__10_), .B(n876), .Y(n1187) );
  OAI221XL U2200 ( .A0(n7330), .A1(n1192), .B0(n51), .B1(n1188), .C0(n1185), 
        .Y(n2153) );
  OAI221XL U2201 ( .A0(n7340), .A1(n1193), .B0(n9290), .B1(n1188), .C0(n1185), 
        .Y(n2121) );
  OAI221XL U2202 ( .A0(n9360), .A1(n1198), .B0(n83), .B1(n1197), .C0(n1196), 
        .Y(n2186) );
  NAND2X1 U2203 ( .A(stg2_real_0__9_), .B(n876), .Y(n1196) );
  OAI221XL U2204 ( .A0(n860), .A1(n1201), .B0(n19), .B1(n1197), .C0(n1194), 
        .Y(n2154) );
  OAI221XL U2205 ( .A0(n859), .A1(n1202), .B0(n9290), .B1(n1197), .C0(n1194), 
        .Y(n2122) );
  OAI221XL U2206 ( .A0(n9370), .A1(n1290), .B0(n76), .B1(n3070), .C0(n1289), 
        .Y(n2244) );
  NAND2X1 U2207 ( .A(stg2_real_2__15_), .B(n880), .Y(n1289) );
  OAI221XL U2208 ( .A0(n9370), .A1(n1295), .B0(n84), .B1(n2710), .C0(n1294), 
        .Y(n2245) );
  NAND2X1 U2209 ( .A(stg2_real_2__14_), .B(n880), .Y(n1294) );
  OAI221XL U2210 ( .A0(n9370), .A1(n1305), .B0(n77), .B1(n1304), .C0(n1303), 
        .Y(n2246) );
  NAND2X1 U2211 ( .A(stg2_real_2__13_), .B(n879), .Y(n1303) );
  OAI221XL U2212 ( .A0(n9370), .A1(n1314), .B0(n81), .B1(n1313), .C0(n1312), 
        .Y(n2247) );
  NAND2X1 U2213 ( .A(stg2_real_2__12_), .B(n879), .Y(n1312) );
  OAI221XL U2214 ( .A0(n9370), .A1(n1323), .B0(n81), .B1(n1322), .C0(n1321), 
        .Y(n2248) );
  NAND2X1 U2215 ( .A(stg2_real_2__11_), .B(n881), .Y(n1321) );
  OAI221XL U2216 ( .A0(n9370), .A1(n1332), .B0(n76), .B1(n1331), .C0(n1330), 
        .Y(n2249) );
  NAND2X1 U2217 ( .A(stg2_real_2__10_), .B(n881), .Y(n1330) );
  OAI221XL U2218 ( .A0(n9370), .A1(n1341), .B0(n79), .B1(n1340), .C0(n1339), 
        .Y(n2250) );
  NAND2X1 U2219 ( .A(stg2_real_2__9_), .B(n881), .Y(n1339) );
  OAI221XL U2220 ( .A0(n9370), .A1(n1350), .B0(n84), .B1(n1349), .C0(n1348), 
        .Y(n2251) );
  NAND2X1 U2221 ( .A(stg2_real_2__8_), .B(n881), .Y(n1348) );
  OAI221XL U2222 ( .A0(n9390), .A1(n2559), .B0(n80), .B1(n2558), .C0(n2557), 
        .Y(n2276) );
  NAND2X1 U2223 ( .A(stg2_real_3__15_), .B(n885), .Y(n2557) );
  OAI221XL U2224 ( .A0(n9400), .A1(n2567), .B0(n83), .B1(n2566), .C0(n2565), 
        .Y(n2277) );
  NAND2X1 U2225 ( .A(stg2_real_3__14_), .B(n884), .Y(n2565) );
  OAI221XL U2226 ( .A0(n9400), .A1(n2576), .B0(n81), .B1(n2575), .C0(n2574), 
        .Y(n2278) );
  NAND2X1 U2227 ( .A(stg2_real_3__13_), .B(n877), .Y(n2574) );
  OAI221XL U2228 ( .A0(n9400), .A1(n2585), .B0(n80), .B1(n2584), .C0(n2583), 
        .Y(n2279) );
  NAND2X1 U2229 ( .A(stg2_real_3__12_), .B(n885), .Y(n2583) );
  OAI221XL U2230 ( .A0(n9400), .A1(n2594), .B0(n81), .B1(n2593), .C0(n2592), 
        .Y(n2280) );
  NAND2X1 U2231 ( .A(stg2_real_3__11_), .B(n884), .Y(n2592) );
  OAI221XL U2232 ( .A0(n9400), .A1(n2603), .B0(n83), .B1(n2602), .C0(n2601), 
        .Y(n2281) );
  NAND2X1 U2233 ( .A(stg2_real_3__10_), .B(n884), .Y(n2601) );
  OAI221XL U2234 ( .A0(n9400), .A1(n2612), .B0(n83), .B1(n2611), .C0(n2610), 
        .Y(n2282) );
  NAND2X1 U2235 ( .A(stg2_real_3__9_), .B(n885), .Y(n2610) );
  OAI221XL U2236 ( .A0(n9400), .A1(n2621), .B0(n78), .B1(n2620), .C0(n2619), 
        .Y(n2283) );
  NAND2X1 U2237 ( .A(stg2_real_3__8_), .B(n884), .Y(n2619) );
  OAI221XL U2238 ( .A0(n9380), .A1(n1426), .B0(n79), .B1(n1425), .C0(n1424), 
        .Y(n2212) );
  NAND2X1 U2239 ( .A(stg2_real_1__15_), .B(n881), .Y(n1424) );
  OAI221XL U2240 ( .A0(n9380), .A1(n1433), .B0(n79), .B1(n1432), .C0(n1431), 
        .Y(n2213) );
  NAND2X1 U2241 ( .A(stg2_real_1__14_), .B(n881), .Y(n1431) );
  OAI221XL U2242 ( .A0(n9380), .A1(n1796), .B0(n78), .B1(n1795), .C0(n1794), 
        .Y(n2214) );
  NAND2X1 U2243 ( .A(stg2_real_1__13_), .B(n883), .Y(n1794) );
  OAI221XL U2244 ( .A0(n9380), .A1(n1803), .B0(n80), .B1(n1802), .C0(n1801), 
        .Y(n2215) );
  NAND2X1 U2245 ( .A(stg2_real_1__12_), .B(n883), .Y(n1801) );
  OAI221XL U2246 ( .A0(n9380), .A1(n1812), .B0(n82), .B1(n1809), .C0(n1808), 
        .Y(n2216) );
  NAND2X1 U2247 ( .A(stg2_real_1__11_), .B(n883), .Y(n1808) );
  OAI221XL U2248 ( .A0(n9390), .A1(n2315), .B0(n78), .B1(n2314), .C0(n2313), 
        .Y(n2217) );
  NAND2X1 U2249 ( .A(stg2_real_1__10_), .B(n883), .Y(n2313) );
  OAI221XL U2250 ( .A0(n9390), .A1(n2322), .B0(n79), .B1(n2321), .C0(n2320), 
        .Y(n2218) );
  NAND2X1 U2251 ( .A(stg2_real_1__9_), .B(n883), .Y(n2320) );
  OAI221XL U2252 ( .A0(n9390), .A1(n2329), .B0(n77), .B1(n2328), .C0(n2327), 
        .Y(n2219) );
  NAND2X1 U2253 ( .A(stg2_real_1__8_), .B(n882), .Y(n2327) );
  CLKINVX1 U2254 ( .A(stg2_img_15__0_), .Y(n3194) );
  CLKINVX1 U2255 ( .A(stg2_img_11__1_), .Y(n3195) );
  CLKINVX1 U2256 ( .A(stg2_img_11__2_), .Y(n3196) );
  CLKINVX1 U2257 ( .A(stg2_img_11__3_), .Y(n3197) );
  CLKINVX1 U2258 ( .A(stg2_img_11__4_), .Y(n3198) );
  CLKINVX1 U2259 ( .A(stg2_img_11__5_), .Y(n3199) );
  CLKINVX1 U2260 ( .A(stg2_img_11__6_), .Y(n3200) );
  CLKINVX1 U2261 ( .A(stg2_img_11__7_), .Y(n3201) );
  CLKINVX1 U2262 ( .A(stg2_img_11__8_), .Y(n3202) );
  CLKINVX1 U2263 ( .A(stg2_img_11__9_), .Y(n3203) );
  CLKINVX1 U2264 ( .A(stg2_img_11__10_), .Y(n3204) );
  CLKINVX1 U2265 ( .A(stg2_img_11__11_), .Y(n3205) );
  CLKINVX1 U2266 ( .A(stg2_img_11__12_), .Y(n3206) );
  OA22X1 U2267 ( .A0(n202), .A1(n2613), .B0(n76), .B1(n2612), .Y(n2614) );
  OA22X1 U2268 ( .A0(n191), .A1(n2604), .B0(n80), .B1(n2603), .Y(n2605) );
  OA22X1 U2269 ( .A0(n189), .A1(n2595), .B0(n80), .B1(n2594), .Y(n2596) );
  OA22X1 U2270 ( .A0(n203), .A1(n2586), .B0(n78), .B1(n2585), .Y(n2587) );
  OA22X1 U2271 ( .A0(n191), .A1(n2577), .B0(n76), .B1(n2576), .Y(n2578) );
  OA22X1 U2272 ( .A0(n189), .A1(n2568), .B0(n83), .B1(n2567), .Y(n2569) );
  OA22X1 U2273 ( .A0(n200), .A1(n2560), .B0(n82), .B1(n2559), .Y(n2561) );
  OA22X1 U2274 ( .A0(n191), .A1(n1351), .B0(n79), .B1(n1350), .Y(n1352) );
  OA22X1 U2275 ( .A0(n205), .A1(n1342), .B0(n75), .B1(n1341), .Y(n1343) );
  OA22X1 U2276 ( .A0(n181), .A1(n1333), .B0(n84), .B1(n1332), .Y(n1334) );
  OA22X1 U2277 ( .A0(n195), .A1(n1324), .B0(n81), .B1(n1323), .Y(n1325) );
  OA22X1 U2278 ( .A0(n183), .A1(n1315), .B0(n80), .B1(n1314), .Y(n1316) );
  OA22X1 U2279 ( .A0(n207), .A1(n1306), .B0(n79), .B1(n1305), .Y(n1307) );
  OA22X1 U2280 ( .A0(n197), .A1(n2708), .B0(n76), .B1(n1295), .Y(n1296) );
  OA22X1 U2281 ( .A0(n205), .A1(n3068), .B0(n75), .B1(n1290), .Y(n1291) );
  OA22X1 U2282 ( .A0(n200), .A1(n1217), .B0(n82), .B1(n1216), .Y(n1218) );
  OA22X1 U2283 ( .A0(n200), .A1(n1208), .B0(n80), .B1(n1207), .Y(n1209) );
  OA22X1 U2284 ( .A0(n205), .A1(n1199), .B0(n78), .B1(n1198), .Y(n1200) );
  OA22X1 U2285 ( .A0(n200), .A1(n1190), .B0(n77), .B1(n1189), .Y(n1191) );
  OA22X1 U2286 ( .A0(n189), .A1(n1181), .B0(n75), .B1(n1180), .Y(n1182) );
  OA22X1 U2287 ( .A0(n185), .A1(n1172), .B0(n82), .B1(n1171), .Y(n1173) );
  OA22X1 U2288 ( .A0(n195), .A1(n1163), .B0(n82), .B1(n1162), .Y(n1164) );
  OA22X1 U2289 ( .A0(n203), .A1(n1154), .B0(n78), .B1(n1153), .Y(n1155) );
  OA22X1 U2290 ( .A0(n199), .A1(n2766), .B0(n81), .B1(n2322), .Y(n2323) );
  OA22X1 U2291 ( .A0(n9630), .A1(n2756), .B0(n79), .B1(n2315), .Y(n2316) );
  OA22X1 U2292 ( .A0(n183), .A1(n2746), .B0(n76), .B1(n1812), .Y(n2309) );
  OA22X1 U2293 ( .A0(n207), .A1(n2736), .B0(n76), .B1(n1803), .Y(n1804) );
  OA22X1 U2294 ( .A0(n187), .A1(n2726), .B0(n84), .B1(n1796), .Y(n1797) );
  OA22X1 U2295 ( .A0(n203), .A1(n2716), .B0(n80), .B1(n1433), .Y(n1434) );
  OA22X1 U2296 ( .A0(n207), .A1(n3074), .B0(n83), .B1(n1426), .Y(n1427) );
  OAI222XL U2297 ( .A0(n897), .A1(n3158), .B0(n860), .B1(n10980), .C0(n47), 
        .C1(n10940), .Y(n2171) );
  OAI222XL U2298 ( .A0(n148), .A1(n898), .B0(n859), .B1(n10990), .C0(n9300), 
        .C1(n10940), .Y(n2139) );
  OAI222XL U2299 ( .A0(n897), .A1(n3157), .B0(n860), .B1(n11040), .C0(n49), 
        .C1(n11000), .Y(n2172) );
  OAI222XL U2300 ( .A0(n149), .A1(n897), .B0(n859), .B1(n11050), .C0(n9300), 
        .C1(n11000), .Y(n2140) );
  OAI222XL U2301 ( .A0(n897), .A1(n3156), .B0(n860), .B1(n11100), .C0(n50), 
        .C1(n11060), .Y(n2173) );
  OAI222XL U2302 ( .A0(n162), .A1(n896), .B0(n859), .B1(n11110), .C0(n9290), 
        .C1(n11060), .Y(n2141) );
  OAI222XL U2303 ( .A0(n897), .A1(n3155), .B0(n860), .B1(n11160), .C0(n20), 
        .C1(n11120), .Y(n2174) );
  OAI222XL U2304 ( .A0(n163), .A1(n895), .B0(n859), .B1(n11170), .C0(n9300), 
        .C1(n11120), .Y(n2142) );
  OAI222XL U2305 ( .A0(n896), .A1(n3154), .B0(n860), .B1(n11220), .C0(n19), 
        .C1(n11180), .Y(n2175) );
  OAI222XL U2306 ( .A0(n164), .A1(n888), .B0(n859), .B1(n11230), .C0(n9320), 
        .C1(n11180), .Y(n2143) );
  OAI222XL U2307 ( .A0(n896), .A1(n3153), .B0(n860), .B1(n11280), .C0(n46), 
        .C1(n11240), .Y(n2176) );
  OAI222XL U2308 ( .A0(n173), .A1(n888), .B0(n859), .B1(n11290), .C0(n9300), 
        .C1(n11240), .Y(n2144) );
  OAI222XL U2309 ( .A0(n896), .A1(n3152), .B0(n860), .B1(n11340), .C0(n47), 
        .C1(n11300), .Y(n2177) );
  OAI222XL U2310 ( .A0(n174), .A1(n888), .B0(n859), .B1(n11350), .C0(n9310), 
        .C1(n11300), .Y(n2145) );
  OAI222XL U2311 ( .A0(n896), .A1(n3151), .B0(n860), .B1(n11400), .C0(n51), 
        .C1(n11360), .Y(n2178) );
  OAI222XL U2312 ( .A0(n172), .A1(n888), .B0(n859), .B1(n11410), .C0(n9300), 
        .C1(n11360), .Y(n2146) );
  OAI222XL U2313 ( .A0(n896), .A1(n3150), .B0(n860), .B1(n1146), .C0(n48), 
        .C1(n11420), .Y(n2179) );
  OAI222XL U2314 ( .A0(n3150), .A1(n898), .B0(n859), .B1(n1147), .C0(n9350), 
        .C1(n11420), .Y(n2147) );
  OAI221XL U2315 ( .A0(n844), .A1(n1280), .B0(n181), .B1(n1278), .C0(n1276), 
        .Y(n3224) );
  NAND2X1 U2316 ( .A(stg2_real_4__0_), .B(n880), .Y(n1276) );
  OAI221XL U2317 ( .A0(n844), .A1(n1217), .B0(n189), .B1(n1215), .C0(n1213), 
        .Y(n3217) );
  NAND2X1 U2318 ( .A(stg2_real_4__7_), .B(n876), .Y(n1213) );
  OAI221XL U2319 ( .A0(n844), .A1(n1226), .B0(n207), .B1(n1224), .C0(n1222), 
        .Y(n3218) );
  NAND2X1 U2320 ( .A(stg2_real_4__6_), .B(n877), .Y(n1222) );
  OAI221XL U2321 ( .A0(n844), .A1(n1235), .B0(n187), .B1(n1233), .C0(n1231), 
        .Y(n3219) );
  NAND2X1 U2322 ( .A(stg2_real_4__5_), .B(n879), .Y(n1231) );
  OAI221XL U2323 ( .A0(n844), .A1(n1244), .B0(n191), .B1(n1242), .C0(n1240), 
        .Y(n3220) );
  NAND2X1 U2324 ( .A(stg2_real_4__4_), .B(n879), .Y(n1240) );
  OAI221XL U2325 ( .A0(n844), .A1(n1253), .B0(n205), .B1(n1251), .C0(n1249), 
        .Y(n3221) );
  NAND2X1 U2326 ( .A(stg2_real_4__3_), .B(n879), .Y(n1249) );
  OAI221XL U2327 ( .A0(n844), .A1(n1262), .B0(n195), .B1(n1260), .C0(n1258), 
        .Y(n3222) );
  NAND2X1 U2328 ( .A(stg2_real_4__2_), .B(n878), .Y(n1258) );
  OAI221XL U2329 ( .A0(n844), .A1(n1271), .B0(n197), .B1(n1269), .C0(n1267), 
        .Y(n3223) );
  NAND2X1 U2330 ( .A(stg2_real_4__1_), .B(n878), .Y(n1267) );
  OAI221XL U2331 ( .A0(n9370), .A1(n1279), .B0(n80), .B1(n1278), .C0(n1277), 
        .Y(n2195) );
  NAND2X1 U2332 ( .A(stg2_real_0__0_), .B(n880), .Y(n1277) );
  OAI221XL U2333 ( .A0(n7330), .A1(n1282), .B0(n20), .B1(n1278), .C0(n1275), 
        .Y(n2163) );
  OAI221XL U2334 ( .A0(n859), .A1(n1283), .B0(n9320), .B1(n1278), .C0(n1275), 
        .Y(n2131) );
  OAI221XL U2335 ( .A0(n9380), .A1(n1414), .B0(n83), .B1(n1413), .C0(n1412), 
        .Y(n2259) );
  NAND2X1 U2336 ( .A(stg2_real_2__0_), .B(n881), .Y(n1412) );
  OAI221XL U2337 ( .A0(n9380), .A1(n2695), .B0(n75), .B1(n2694), .C0(n2693), 
        .Y(n2291) );
  NAND2X1 U2338 ( .A(stg2_real_3__0_), .B(n886), .Y(n2693) );
  OAI221XL U2339 ( .A0(n9390), .A1(n2385), .B0(n84), .B1(n2384), .C0(n2383), 
        .Y(n2227) );
  NAND2X1 U2340 ( .A(stg2_real_1__0_), .B(n886), .Y(n2383) );
  OAI221XL U2341 ( .A0(n9360), .A1(n1207), .B0(n75), .B1(n1206), .C0(n1205), 
        .Y(n2187) );
  NAND2X1 U2342 ( .A(stg2_real_0__8_), .B(n876), .Y(n1205) );
  OAI221XL U2343 ( .A0(n860), .A1(n1210), .B0(n50), .B1(n1206), .C0(n1203), 
        .Y(n2155) );
  OAI221XL U2344 ( .A0(n859), .A1(n1211), .B0(n9310), .B1(n1206), .C0(n1203), 
        .Y(n2123) );
  OAI221XL U2345 ( .A0(n9360), .A1(n1216), .B0(n81), .B1(n1215), .C0(n1214), 
        .Y(n2188) );
  NAND2X1 U2346 ( .A(stg2_real_0__7_), .B(n876), .Y(n1214) );
  OAI221XL U2347 ( .A0(n860), .A1(n1219), .B0(n50), .B1(n1215), .C0(n1212), 
        .Y(n2156) );
  OAI221XL U2348 ( .A0(n859), .A1(n1220), .B0(n9330), .B1(n1215), .C0(n1212), 
        .Y(n2124) );
  OAI221XL U2349 ( .A0(n9360), .A1(n1225), .B0(n81), .B1(n1224), .C0(n1223), 
        .Y(n2189) );
  NAND2X1 U2350 ( .A(stg2_real_0__6_), .B(n877), .Y(n1223) );
  OAI221XL U2351 ( .A0(n7330), .A1(n1228), .B0(n52), .B1(n1224), .C0(n1221), 
        .Y(n2157) );
  OAI221XL U2352 ( .A0(n859), .A1(n1229), .B0(n9350), .B1(n1224), .C0(n1221), 
        .Y(n2125) );
  OAI221XL U2353 ( .A0(n9360), .A1(n1234), .B0(n80), .B1(n1233), .C0(n1232), 
        .Y(n2190) );
  NAND2X1 U2354 ( .A(stg2_real_0__5_), .B(n879), .Y(n1232) );
  OAI221XL U2355 ( .A0(n7330), .A1(n1237), .B0(n48), .B1(n1233), .C0(n1230), 
        .Y(n2158) );
  OAI221XL U2356 ( .A0(n859), .A1(n1238), .B0(n9350), .B1(n1233), .C0(n1230), 
        .Y(n2126) );
  OAI221XL U2357 ( .A0(n9360), .A1(n1243), .B0(n82), .B1(n1242), .C0(n1241), 
        .Y(n2191) );
  NAND2X1 U2358 ( .A(stg2_real_0__4_), .B(n879), .Y(n1241) );
  OAI221XL U2359 ( .A0(n860), .A1(n1246), .B0(n20), .B1(n1242), .C0(n1239), 
        .Y(n2159) );
  OAI221XL U2360 ( .A0(n859), .A1(n1247), .B0(n9340), .B1(n1242), .C0(n1239), 
        .Y(n2127) );
  OAI221XL U2361 ( .A0(n9360), .A1(n1252), .B0(n78), .B1(n1251), .C0(n1250), 
        .Y(n2192) );
  NAND2X1 U2362 ( .A(stg2_real_0__3_), .B(n878), .Y(n1250) );
  OAI221XL U2363 ( .A0(n860), .A1(n1255), .B0(n52), .B1(n1251), .C0(n1248), 
        .Y(n2160) );
  OAI221XL U2364 ( .A0(n7340), .A1(n1256), .B0(n9350), .B1(n1251), .C0(n1248), 
        .Y(n2128) );
  OAI221XL U2365 ( .A0(n9370), .A1(n1261), .B0(n76), .B1(n1260), .C0(n1259), 
        .Y(n2193) );
  NAND2X1 U2366 ( .A(stg2_real_0__2_), .B(n882), .Y(n1259) );
  OAI221XL U2367 ( .A0(n860), .A1(n1264), .B0(n20), .B1(n1260), .C0(n1257), 
        .Y(n2161) );
  OAI221XL U2368 ( .A0(n7340), .A1(n1265), .B0(n9350), .B1(n1260), .C0(n1257), 
        .Y(n2129) );
  OAI221XL U2369 ( .A0(n9370), .A1(n1270), .B0(n75), .B1(n1269), .C0(n1268), 
        .Y(n2194) );
  NAND2X1 U2370 ( .A(stg2_real_0__1_), .B(n880), .Y(n1268) );
  OAI221XL U2371 ( .A0(n860), .A1(n1273), .B0(n50), .B1(n1269), .C0(n1266), 
        .Y(n2162) );
  OAI221XL U2372 ( .A0(n7340), .A1(n1274), .B0(n9330), .B1(n1269), .C0(n1266), 
        .Y(n2130) );
  OAI221XL U2373 ( .A0(n9370), .A1(n1358), .B0(n76), .B1(n1357), .C0(n1356), 
        .Y(n2252) );
  NAND2X1 U2374 ( .A(stg2_real_2__7_), .B(n880), .Y(n1356) );
  OAI221XL U2375 ( .A0(n9380), .A1(n1366), .B0(n83), .B1(n1365), .C0(n1364), 
        .Y(n2253) );
  NAND2X1 U2376 ( .A(stg2_real_2__6_), .B(n880), .Y(n1364) );
  OAI221XL U2377 ( .A0(n9380), .A1(n1374), .B0(n76), .B1(n1373), .C0(n1372), 
        .Y(n2254) );
  NAND2X1 U2378 ( .A(stg2_real_2__5_), .B(n880), .Y(n1372) );
  OAI221XL U2379 ( .A0(n9380), .A1(n1382), .B0(n77), .B1(n1381), .C0(n1380), 
        .Y(n2255) );
  NAND2X1 U2380 ( .A(stg2_real_2__4_), .B(n882), .Y(n1380) );
  OAI221XL U2381 ( .A0(n9380), .A1(n1390), .B0(n78), .B1(n1389), .C0(n1388), 
        .Y(n2256) );
  NAND2X1 U2382 ( .A(stg2_real_2__3_), .B(n882), .Y(n1388) );
  OAI221XL U2383 ( .A0(n9380), .A1(n1398), .B0(n78), .B1(n1397), .C0(n1396), 
        .Y(n2257) );
  NAND2X1 U2384 ( .A(stg2_real_2__2_), .B(n882), .Y(n1396) );
  OAI221XL U2385 ( .A0(n9380), .A1(n1406), .B0(n77), .B1(n1405), .C0(n1404), 
        .Y(n2258) );
  NAND2X1 U2386 ( .A(stg2_real_2__1_), .B(n882), .Y(n1404) );
  OAI221XL U2387 ( .A0(n9400), .A1(n2630), .B0(n75), .B1(n2629), .C0(n2628), 
        .Y(n2284) );
  NAND2X1 U2388 ( .A(stg2_real_3__7_), .B(n885), .Y(n2628) );
  OAI221XL U2389 ( .A0(n9400), .A1(n2639), .B0(n84), .B1(n2638), .C0(n2637), 
        .Y(n2285) );
  NAND2X1 U2390 ( .A(stg2_real_3__6_), .B(n886), .Y(n2637) );
  OAI221XL U2391 ( .A0(n9400), .A1(n2648), .B0(n84), .B1(n2647), .C0(n2646), 
        .Y(n2286) );
  NAND2X1 U2392 ( .A(stg2_real_3__5_), .B(n878), .Y(n2646) );
  OAI221XL U2393 ( .A0(n9400), .A1(n2657), .B0(n83), .B1(n2656), .C0(n2655), 
        .Y(n2287) );
  NAND2X1 U2394 ( .A(stg2_real_3__4_), .B(n885), .Y(n2655) );
  OAI221XL U2395 ( .A0(n9400), .A1(n2666), .B0(n79), .B1(n2665), .C0(n2664), 
        .Y(n2288) );
  NAND2X1 U2396 ( .A(stg2_real_3__3_), .B(n878), .Y(n2664) );
  OAI221XL U2397 ( .A0(n9380), .A1(n2675), .B0(n84), .B1(n2674), .C0(n2673), 
        .Y(n2289) );
  NAND2X1 U2398 ( .A(stg2_real_3__2_), .B(n885), .Y(n2673) );
  OAI221XL U2399 ( .A0(n9380), .A1(n2684), .B0(n79), .B1(n2683), .C0(n2682), 
        .Y(n2290) );
  NAND2X1 U2400 ( .A(stg2_real_3__1_), .B(n885), .Y(n2682) );
  OAI221XL U2401 ( .A0(n9390), .A1(n2336), .B0(n81), .B1(n2335), .C0(n2334), 
        .Y(n2220) );
  NAND2X1 U2402 ( .A(stg2_real_1__7_), .B(n882), .Y(n2334) );
  OAI221XL U2403 ( .A0(n9390), .A1(n2343), .B0(n82), .B1(n2342), .C0(n2341), 
        .Y(n2221) );
  NAND2X1 U2404 ( .A(stg2_real_1__6_), .B(n884), .Y(n2341) );
  OAI221XL U2405 ( .A0(n9390), .A1(n2350), .B0(n82), .B1(n2349), .C0(n2348), 
        .Y(n2222) );
  NAND2X1 U2406 ( .A(stg2_real_1__5_), .B(n884), .Y(n2348) );
  OAI221XL U2407 ( .A0(n9390), .A1(n2357), .B0(n76), .B1(n2356), .C0(n2355), 
        .Y(n2223) );
  NAND2X1 U2408 ( .A(stg2_real_1__4_), .B(n884), .Y(n2355) );
  OAI221XL U2409 ( .A0(n9390), .A1(n2364), .B0(n80), .B1(n2363), .C0(n2362), 
        .Y(n2224) );
  NAND2X1 U2410 ( .A(stg2_real_1__3_), .B(n883), .Y(n2362) );
  OAI221XL U2411 ( .A0(n9390), .A1(n2371), .B0(n78), .B1(n2370), .C0(n2369), 
        .Y(n2225) );
  NAND2X1 U2412 ( .A(stg2_real_1__2_), .B(n883), .Y(n2369) );
  OAI221XL U2413 ( .A0(n9390), .A1(n2378), .B0(n82), .B1(n2377), .C0(n2376), 
        .Y(n2226) );
  NAND2X1 U2414 ( .A(stg2_real_1__1_), .B(n877), .Y(n2376) );
  CLKINVX1 U2415 ( .A(stg2_img_11__13_), .Y(n3207) );
  CLKINVX1 U2416 ( .A(stg2_img_11__14_), .Y(n3208) );
  OA22X1 U2417 ( .A0(n199), .A1(n2704), .B0(n76), .B1(n2703), .Y(n2705) );
  NAND2X1 U2418 ( .A(stg2_real_12__14_), .B(n877), .Y(n1148) );
  NAND2X1 U2419 ( .A(stg2_real_12__13_), .B(n877), .Y(n1158) );
  NAND2X1 U2420 ( .A(stg2_real_12__12_), .B(n877), .Y(n1167) );
  NAND2X1 U2421 ( .A(stg2_real_12__11_), .B(n878), .Y(n1176) );
  NAND2X1 U2422 ( .A(stg2_real_12__10_), .B(n878), .Y(n1185) );
  AND2X2 U2423 ( .A(stg2_img_15__0_), .B(n885), .Y(n792) );
  CLKINVX1 U2424 ( .A(stg2_img_8__0_), .Y(n3150) );
  AND2X2 U2425 ( .A(stg2_img_14__0_), .B(n886), .Y(n793) );
  AND2X2 U2426 ( .A(stg2_real_13__14_), .B(n881), .Y(n794) );
  AND2X2 U2427 ( .A(stg2_real_13__13_), .B(n881), .Y(n795) );
  AND2X2 U2428 ( .A(stg2_real_13__12_), .B(n883), .Y(n796) );
  AND2X2 U2429 ( .A(stg2_real_13__11_), .B(n883), .Y(n797) );
  AND2X2 U2430 ( .A(stg2_real_13__10_), .B(n883), .Y(n798) );
  AND2X2 U2431 ( .A(stg2_real_13__9_), .B(n883), .Y(n799) );
  AND2X2 U2432 ( .A(stg2_real_13__8_), .B(n882), .Y(n800) );
  AND2X2 U2433 ( .A(stg2_real_13__7_), .B(n882), .Y(n801) );
  AND2X2 U2434 ( .A(stg2_real_13__6_), .B(n882), .Y(n802) );
  AND2X2 U2435 ( .A(stg2_real_13__5_), .B(n884), .Y(n803) );
  AND2X2 U2436 ( .A(stg2_real_13__4_), .B(n884), .Y(n804) );
  AND2X2 U2437 ( .A(stg2_real_13__3_), .B(n883), .Y(n805) );
  AND2X2 U2438 ( .A(stg2_real_13__2_), .B(n883), .Y(n806) );
  AND2X2 U2439 ( .A(stg2_real_13__1_), .B(n883), .Y(n807) );
  AND2X2 U2440 ( .A(stg2_real_14__14_), .B(n880), .Y(n808) );
  AND2X2 U2441 ( .A(stg2_real_14__13_), .B(n879), .Y(n809) );
  AND2X2 U2442 ( .A(stg2_real_14__12_), .B(n879), .Y(n810) );
  AND2X2 U2443 ( .A(stg2_real_14__11_), .B(n879), .Y(n811) );
  AND2X2 U2444 ( .A(stg2_real_14__10_), .B(n881), .Y(n812) );
  AND2X2 U2445 ( .A(stg2_real_14__9_), .B(n881), .Y(n813) );
  AND2X2 U2446 ( .A(stg2_real_14__8_), .B(n881), .Y(n814) );
  AND2X2 U2447 ( .A(stg2_real_14__7_), .B(n881), .Y(n815) );
  AND2X2 U2448 ( .A(stg2_real_14__6_), .B(n880), .Y(n816) );
  AND2X2 U2449 ( .A(stg2_real_14__5_), .B(n880), .Y(n817) );
  AND2X2 U2450 ( .A(stg2_real_14__4_), .B(n880), .Y(n818) );
  AND2X2 U2451 ( .A(stg2_real_14__3_), .B(n882), .Y(n819) );
  AND2X2 U2452 ( .A(stg2_real_14__2_), .B(n882), .Y(n820) );
  AND2X2 U2453 ( .A(stg2_real_14__1_), .B(n882), .Y(n821) );
  AND2X2 U2454 ( .A(stg2_real_15__14_), .B(n884), .Y(n822) );
  AND2X2 U2455 ( .A(stg2_real_15__10_), .B(n884), .Y(n823) );
  AND2X2 U2456 ( .A(stg2_real_15__9_), .B(n884), .Y(n824) );
  AND2X2 U2457 ( .A(stg2_real_15__8_), .B(n884), .Y(n825) );
  AND2X2 U2458 ( .A(stg2_real_15__7_), .B(n878), .Y(n826) );
  AND2X2 U2459 ( .A(stg2_real_15__6_), .B(n886), .Y(n827) );
  AND2X2 U2460 ( .A(stg2_real_15__5_), .B(n878), .Y(n828) );
  AND2X2 U2461 ( .A(stg2_real_15__4_), .B(n886), .Y(n829) );
  AND2X2 U2462 ( .A(stg2_real_15__3_), .B(n886), .Y(n830) );
  AND2X2 U2463 ( .A(stg2_img_13__0_), .B(n878), .Y(n831) );
  CLKINVX1 U2464 ( .A(stg2_img_14__0_), .Y(n3181) );
  CLKINVX1 U2465 ( .A(stg2_img_13__0_), .Y(n3166) );
  AND2X2 U2466 ( .A(stg2_real_15__13_), .B(n885), .Y(n832) );
  AND2X2 U2467 ( .A(stg2_real_15__12_), .B(n885), .Y(n833) );
  AND2X2 U2468 ( .A(stg2_real_15__11_), .B(n885), .Y(n834) );
  AND2X2 U2469 ( .A(stg2_real_15__2_), .B(n885), .Y(n835) );
  AND2X2 U2470 ( .A(stg2_real_15__1_), .B(n885), .Y(n836) );
  CLKINVX1 U2471 ( .A(stg2_img_8__1_), .Y(n3151) );
  CLKINVX1 U2472 ( .A(stg2_img_10__1_), .Y(n3182) );
  CLKINVX1 U2473 ( .A(stg2_img_9__1_), .Y(n3167) );
  CLKINVX1 U2474 ( .A(stg2_img_8__2_), .Y(n3152) );
  CLKINVX1 U2475 ( .A(stg2_img_10__2_), .Y(n3183) );
  CLKINVX1 U2476 ( .A(stg2_img_9__2_), .Y(n3168) );
  CLKINVX1 U2477 ( .A(stg2_img_8__3_), .Y(n3153) );
  CLKINVX1 U2478 ( .A(stg2_img_10__3_), .Y(n3184) );
  CLKINVX1 U2479 ( .A(stg2_img_9__3_), .Y(n3169) );
  CLKINVX1 U2480 ( .A(stg2_img_8__4_), .Y(n3154) );
  CLKINVX1 U2481 ( .A(stg2_img_10__4_), .Y(n3185) );
  CLKINVX1 U2482 ( .A(stg2_img_9__4_), .Y(n3170) );
  CLKINVX1 U2483 ( .A(stg2_img_8__5_), .Y(n3155) );
  CLKINVX1 U2484 ( .A(stg2_img_10__5_), .Y(n3186) );
  CLKINVX1 U2485 ( .A(stg2_img_9__5_), .Y(n3171) );
  CLKINVX1 U2486 ( .A(stg2_img_8__6_), .Y(n3156) );
  CLKINVX1 U2487 ( .A(stg2_img_10__6_), .Y(n3187) );
  CLKINVX1 U2488 ( .A(stg2_img_9__6_), .Y(n3172) );
  CLKINVX1 U2489 ( .A(stg2_img_8__7_), .Y(n3157) );
  CLKINVX1 U2490 ( .A(stg2_img_10__7_), .Y(n3188) );
  CLKINVX1 U2491 ( .A(stg2_img_9__7_), .Y(n3173) );
  CLKINVX1 U2492 ( .A(stg2_img_8__8_), .Y(n3158) );
  CLKINVX1 U2493 ( .A(stg2_img_10__8_), .Y(n3189) );
  CLKINVX1 U2494 ( .A(stg2_img_9__8_), .Y(n3174) );
  CLKINVX1 U2495 ( .A(stg2_img_8__9_), .Y(n3159) );
  CLKINVX1 U2496 ( .A(stg2_img_10__9_), .Y(n3190) );
  CLKINVX1 U2497 ( .A(stg2_img_9__9_), .Y(n3175) );
  CLKINVX1 U2498 ( .A(stg2_img_8__10_), .Y(n3160) );
  CLKINVX1 U2499 ( .A(stg2_img_10__10_), .Y(n3191) );
  CLKINVX1 U2500 ( .A(stg2_img_9__10_), .Y(n3176) );
  CLKINVX1 U2501 ( .A(stg2_img_8__11_), .Y(n3161) );
  CLKINVX1 U2502 ( .A(stg2_img_10__11_), .Y(n3192) );
  CLKINVX1 U2503 ( .A(stg2_img_9__11_), .Y(n3177) );
  CLKINVX1 U2504 ( .A(stg2_img_8__12_), .Y(n3162) );
  CLKINVX1 U2505 ( .A(stg2_img_10__12_), .Y(n3193) );
  CLKINVX1 U2506 ( .A(stg2_img_9__12_), .Y(n3178) );
  CLKINVX1 U2507 ( .A(stg2_img_8__13_), .Y(n3163) );
  CLKINVX1 U2508 ( .A(stg2_img_9__13_), .Y(n3179) );
  CLKINVX1 U2509 ( .A(stg2_img_8__14_), .Y(n3164) );
  CLKINVX1 U2510 ( .A(stg2_img_9__14_), .Y(n3180) );
  NAND2X1 U2511 ( .A(stg2_real_12__9_), .B(n876), .Y(n1194) );
  NAND2X1 U2512 ( .A(stg2_real_12__8_), .B(n876), .Y(n1203) );
  NAND2X1 U2513 ( .A(stg2_real_12__7_), .B(n876), .Y(n1212) );
  NAND2X1 U2514 ( .A(stg2_real_12__6_), .B(n877), .Y(n1221) );
  NAND2X1 U2515 ( .A(stg2_real_12__5_), .B(n879), .Y(n1230) );
  NAND2X1 U2516 ( .A(stg2_real_12__4_), .B(n879), .Y(n1239) );
  NAND2X1 U2517 ( .A(stg2_real_12__3_), .B(n879), .Y(n1248) );
  NAND2X1 U2518 ( .A(stg2_real_12__2_), .B(n878), .Y(n1257) );
  NAND2X1 U2519 ( .A(stg2_real_12__1_), .B(n877), .Y(n1266) );
  AOI222XL U2520 ( .A0(stg_reg[37]), .A1(n861), .B0(n914), .B1(stg_reg[69]), 
        .C0(n904), .C1(n1567), .Y(n3001) );
  OA22X1 U2521 ( .A0(n80), .A1(n2971), .B0(n10460), .B1(n2970), .Y(n2972) );
  OA22X1 U2522 ( .A0(n3115), .A1(n9280), .B0(n3072), .B1(n2967), .Y(n2974) );
  OA22X1 U2523 ( .A0(n83), .A1(n2945), .B0(n10350), .B1(n2944), .Y(n2946) );
  OA22X1 U2524 ( .A0(n3106), .A1(n9280), .B0(n9210), .B1(n2941), .Y(n2948) );
  OA22X1 U2525 ( .A0(n81), .A1(n2746), .B0(n10460), .B1(n2745), .Y(n2747) );
  OA22X1 U2526 ( .A0(n50), .A1(n2744), .B0(n193), .B1(n2743), .Y(n2748) );
  OA22X1 U2527 ( .A0(n84), .A1(n2726), .B0(n10460), .B1(n2725), .Y(n2727) );
  OA22X1 U2528 ( .A0(n19), .A1(n2724), .B0(n185), .B1(n2723), .Y(n2728) );
  AOI222XL U2529 ( .A0(stg_reg[43]), .A1(n861), .B0(n914), .B1(stg_reg[75]), 
        .C0(n905), .C1(n1540), .Y(n2923) );
  AOI222XL U2530 ( .A0(stg_reg[45]), .A1(n861), .B0(n914), .B1(stg_reg[77]), 
        .C0(n905), .C1(n1546), .Y(n2897) );
  AOI222XL U2531 ( .A0(stg_reg[62]), .A1(n862), .B0(stg_reg[94]), .B1(n913), 
        .C0(n1725), .C1(n904), .Y(n2720) );
  AOI222XL U2532 ( .A0(stg_reg[46]), .A1(n861), .B0(n914), .B1(stg_reg[78]), 
        .C0(n905), .C1(n1549), .Y(n2885) );
  OA22X1 U2533 ( .A0(n78), .A1(n3036), .B0(n10460), .B1(n3035), .Y(n3037) );
  OA22X1 U2534 ( .A0(n3137), .A1(n9280), .B0(n3072), .B1(n3032), .Y(n3039) );
  OA22X1 U2535 ( .A0(n81), .A1(n3010), .B0(n10460), .B1(n3009), .Y(n3011) );
  OA22X1 U2536 ( .A0(n3129), .A1(n9280), .B0(n3072), .B1(n3006), .Y(n3013) );
  OA22X1 U2537 ( .A0(n80), .A1(n2816), .B0(n10460), .B1(n2815), .Y(n2817) );
  OA22X1 U2538 ( .A0(n48), .A1(n2814), .B0(n189), .B1(n2813), .Y(n2818) );
  OA22X1 U2539 ( .A0(n77), .A1(n2836), .B0(n10350), .B1(n2835), .Y(n2837) );
  OA22X1 U2540 ( .A0(n45), .A1(n2834), .B0(n202), .B1(n2833), .Y(n2838) );
  OA22X1 U2541 ( .A0(n82), .A1(n2958), .B0(n10460), .B1(n2957), .Y(n2959) );
  OA22X1 U2542 ( .A0(n19), .A1(n2794), .B0(n191), .B1(n2793), .Y(n2798) );
  OA22X1 U2543 ( .A0(n83), .A1(n2776), .B0(n10460), .B1(n2775), .Y(n2777) );
  OA22X1 U2544 ( .A0(n79), .A1(n2756), .B0(n10460), .B1(n2755), .Y(n2757) );
  OA22X1 U2545 ( .A0(n47), .A1(n2754), .B0(n200), .B1(n2753), .Y(n2758) );
  NAND4X1 U2546 ( .A(n2740), .B(n2739), .C(n2738), .D(n2737), .Y(mul_2_in[12])
         );
  OA22X1 U2547 ( .A0(n76), .A1(n2736), .B0(n10350), .B1(n2735), .Y(n2737) );
  AOI222XL U2548 ( .A0(stg_reg[60]), .A1(n862), .B0(stg_reg[92]), .B1(n913), 
        .C0(n1719), .C1(n904), .Y(n2740) );
  OA22X1 U2549 ( .A0(n46), .A1(n2734), .B0(n183), .B1(n2733), .Y(n2738) );
  NAND4X1 U2550 ( .A(n2936), .B(n2935), .C(n2934), .D(n2933), .Y(mul_1_in[10])
         );
  OA22X1 U2551 ( .A0(n81), .A1(n2932), .B0(n10460), .B1(n2931), .Y(n2933) );
  AOI222XL U2552 ( .A0(stg_reg[42]), .A1(n861), .B0(n914), .B1(stg_reg[74]), 
        .C0(n905), .C1(n1537), .Y(n2936) );
  OA22X1 U2553 ( .A0(n3102), .A1(n9280), .B0(n9210), .B1(n2928), .Y(n2935) );
  NAND4X1 U2554 ( .A(n2910), .B(n2909), .C(n2908), .D(n2907), .Y(mul_1_in[12])
         );
  OA22X1 U2555 ( .A0(n84), .A1(n2906), .B0(n10460), .B1(n2905), .Y(n2907) );
  AOI222XL U2556 ( .A0(stg_reg[44]), .A1(n861), .B0(n914), .B1(stg_reg[76]), 
        .C0(n905), .C1(n1543), .Y(n2910) );
  OA22X1 U2557 ( .A0(n3094), .A1(n9280), .B0(n918), .B1(n2902), .Y(n2909) );
  OA22X1 U2558 ( .A0(n185), .A1(n3063), .B0(n82), .B1(n2462), .Y(n2463) );
  CLKINVX1 U2559 ( .A(stg_reg[31]), .Y(n3073) );
  CLKINVX1 U2560 ( .A(stg_reg[15]), .Y(n2869) );
  CLKINVX1 U2561 ( .A(n1504), .Y(n2868) );
  CLKINVX1 U2562 ( .A(stg_reg[111]), .Y(n2870) );
  CLKINVX1 U2563 ( .A(stg_reg[127]), .Y(n3074) );
  OA22X1 U2564 ( .A0(n200), .A1(n1144), .B0(n80), .B1(n1143), .Y(n1145) );
  CLKINVX1 U2565 ( .A(stg_reg[128]), .Y(n1144) );
  OA22X1 U2566 ( .A0(n207), .A1(n3139), .B0(n83), .B1(n3138), .Y(n3140) );
  OA22X1 U2567 ( .A0(n9590), .A1(n2546), .B0(n80), .B1(n2545), .Y(n2547) );
  OA22X1 U2568 ( .A0(n197), .A1(n2540), .B0(n75), .B1(n2539), .Y(n2541) );
  OA22X1 U2569 ( .A0(n187), .A1(n2534), .B0(n75), .B1(n2533), .Y(n2535) );
  OA22X1 U2570 ( .A0(n207), .A1(n2528), .B0(n81), .B1(n2527), .Y(n2529) );
  OA22X1 U2571 ( .A0(n200), .A1(n2522), .B0(n80), .B1(n2521), .Y(n2523) );
  OA22X1 U2572 ( .A0(n199), .A1(n2516), .B0(n77), .B1(n2515), .Y(n2517) );
  OA22X1 U2573 ( .A0(n185), .A1(n3113), .B0(n79), .B1(n3112), .Y(n3114) );
  OA22X1 U2574 ( .A0(n185), .A1(n2510), .B0(n78), .B1(n2509), .Y(n2511) );
  OA22X1 U2575 ( .A0(n183), .A1(n2504), .B0(n83), .B1(n2503), .Y(n2505) );
  OAI221X1 U2576 ( .A0(n9790), .A1(n3062), .B0(n19), .B1(n3059), .C0(n2553), 
        .Y(stg2_img_Wn[0]) );
  OA22X1 U2577 ( .A0(n200), .A1(n2552), .B0(n81), .B1(n2551), .Y(n2553) );
  OAI221X1 U2578 ( .A0(n9760), .A1(n3147), .B0(n51), .B1(n114), .C0(n3146), 
        .Y(stg2_img_Wn[16]) );
  OA22X1 U2579 ( .A0(n203), .A1(n3145), .B0(n79), .B1(n3143), .Y(n3146) );
  OA22X1 U2580 ( .A0(n207), .A1(n3049), .B0(n76), .B1(n2454), .Y(n2455) );
  OA22X1 U2581 ( .A0(n191), .A1(n11380), .B0(n83), .B1(n11370), .Y(n11390) );
  CLKINVX1 U2582 ( .A(stg_reg[129]), .Y(n11380) );
  OA22X1 U2583 ( .A0(n205), .A1(n3036), .B0(n79), .B1(n2449), .Y(n2450) );
  OA22X1 U2584 ( .A0(n187), .A1(n11320), .B0(n81), .B1(n11310), .Y(n11330) );
  CLKINVX1 U2585 ( .A(stg_reg[130]), .Y(n11320) );
  OA22X1 U2586 ( .A0(n207), .A1(n3023), .B0(n78), .B1(n2444), .Y(n2445) );
  OA22X1 U2587 ( .A0(n203), .A1(n11260), .B0(n79), .B1(n11250), .Y(n11270) );
  CLKINVX1 U2588 ( .A(stg_reg[131]), .Y(n11260) );
  OA22X1 U2589 ( .A0(n195), .A1(n11200), .B0(n77), .B1(n11190), .Y(n11210) );
  CLKINVX1 U2590 ( .A(stg_reg[132]), .Y(n11200) );
  OA22X1 U2591 ( .A0(n191), .A1(n11140), .B0(n75), .B1(n11130), .Y(n11150) );
  CLKINVX1 U2592 ( .A(stg_reg[133]), .Y(n11140) );
  OA22X1 U2593 ( .A0(n205), .A1(n11080), .B0(n83), .B1(n11070), .Y(n11090) );
  CLKINVX1 U2594 ( .A(stg_reg[134]), .Y(n11080) );
  OA22X1 U2595 ( .A0(n197), .A1(n11020), .B0(n81), .B1(n11010), .Y(n11030) );
  CLKINVX1 U2596 ( .A(stg_reg[135]), .Y(n11020) );
  AO22X1 U2597 ( .A0(n1578), .A1(n9460), .B0(stg4_img[25]), .B1(n60), .Y(n2266) );
  AO22X1 U2598 ( .A0(n1593), .A1(n9440), .B0(stg4_img[15]), .B1(n56), .Y(n2292) );
  AO22X1 U2599 ( .A0(n1591), .A1(n9430), .B0(stg4_img[14]), .B1(n70), .Y(n2293) );
  AO22X1 U2600 ( .A0(n1589), .A1(n9440), .B0(stg4_img[13]), .B1(n64), .Y(n2294) );
  AO22X1 U2601 ( .A0(n1587), .A1(n9440), .B0(stg4_img[12]), .B1(n60), .Y(n2295) );
  AO22X1 U2602 ( .A0(n1585), .A1(n9440), .B0(stg4_img[11]), .B1(n58), .Y(n2296) );
  AO22X1 U2603 ( .A0(n1583), .A1(n9440), .B0(stg4_img[10]), .B1(n70), .Y(n2297) );
  AO22X1 U2604 ( .A0(n1611), .A1(n9440), .B0(stg4_img[9]), .B1(n56), .Y(n2298)
         );
  AO22X1 U2605 ( .A0(n1551), .A1(n9460), .B0(stg4_img[31]), .B1(n72), .Y(n2260) );
  AO22X1 U2606 ( .A0(n1548), .A1(n9460), .B0(stg4_img[30]), .B1(n58), .Y(n2261) );
  AO22X1 U2607 ( .A0(n1545), .A1(n9460), .B0(stg4_img[29]), .B1(n54), .Y(n2262) );
  AO22X1 U2608 ( .A0(n1542), .A1(n9460), .B0(stg4_img[28]), .B1(n68), .Y(n2263) );
  AO22X1 U2609 ( .A0(n1539), .A1(n9460), .B0(stg4_img[27]), .B1(n60), .Y(n2264) );
  AO22X1 U2610 ( .A0(n1536), .A1(n9460), .B0(stg4_img[26]), .B1(n68), .Y(n2265) );
  AO22X1 U2611 ( .A0(n1503), .A1(n9420), .B0(stg4_img[47]), .B1(n62), .Y(n2228) );
  AO22X1 U2612 ( .A0(n1500), .A1(n9420), .B0(stg4_img[46]), .B1(n58), .Y(n2229) );
  AO22X1 U2613 ( .A0(n1497), .A1(n9430), .B0(stg4_img[45]), .B1(n60), .Y(n2230) );
  AO22X1 U2614 ( .A0(n1494), .A1(n9430), .B0(stg4_img[44]), .B1(n64), .Y(n2231) );
  AO22X1 U2615 ( .A0(n1491), .A1(n9430), .B0(stg4_img[43]), .B1(n56), .Y(n2232) );
  AO22X1 U2616 ( .A0(n1488), .A1(n9430), .B0(stg4_img[42]), .B1(n54), .Y(n2233) );
  AO22X1 U2617 ( .A0(n1530), .A1(n9430), .B0(stg4_img[41]), .B1(n54), .Y(n2234) );
  AO22X1 U2618 ( .A0(n1455), .A1(n9420), .B0(stg4_img[63]), .B1(n58), .Y(n2196) );
  AO22X1 U2619 ( .A0(n1452), .A1(n9410), .B0(stg4_img[62]), .B1(n60), .Y(n2197) );
  AO22X1 U2620 ( .A0(n1449), .A1(n9410), .B0(stg4_img[61]), .B1(n66), .Y(n2198) );
  AO22X1 U2621 ( .A0(n1440), .A1(n9450), .B0(stg4_img[58]), .B1(n62), .Y(n2201) );
  AO22X1 U2622 ( .A0(n1482), .A1(n9410), .B0(stg4_img[57]), .B1(n70), .Y(n2202) );
  OA22X1 U2623 ( .A0(n202), .A1(n3103), .B0(n83), .B1(n127), .Y(n3104) );
  OA22X1 U2624 ( .A0(n189), .A1(n2498), .B0(n82), .B1(n128), .Y(n2499) );
  OA22X1 U2625 ( .A0(n195), .A1(n3099), .B0(n83), .B1(n133), .Y(n3100) );
  OA22X1 U2626 ( .A0(n191), .A1(n2493), .B0(n82), .B1(n134), .Y(n2494) );
  OA22X1 U2627 ( .A0(n187), .A1(n3095), .B0(n79), .B1(n135), .Y(n3096) );
  OA22X1 U2628 ( .A0(n185), .A1(n2488), .B0(n78), .B1(n136), .Y(n2489) );
  OA22X1 U2629 ( .A0(n202), .A1(n3091), .B0(n77), .B1(n137), .Y(n3092) );
  OA22X1 U2630 ( .A0(n197), .A1(n2483), .B0(n84), .B1(n138), .Y(n2484) );
  OA22X1 U2631 ( .A0(n193), .A1(n3088), .B0(n75), .B1(n154), .Y(n3089) );
  OA22X1 U2632 ( .A0(n187), .A1(n2478), .B0(n83), .B1(n155), .Y(n2479) );
  OA22X1 U2633 ( .A0(n181), .A1(n3086), .B0(n77), .B1(n156), .Y(n3087) );
  OA22X1 U2634 ( .A0(n199), .A1(n2473), .B0(n81), .B1(n157), .Y(n2474) );
  OA22X1 U2635 ( .A0(n202), .A1(n3084), .B0(n79), .B1(n168), .Y(n3085) );
  OA22X1 U2636 ( .A0(n183), .A1(n2468), .B0(n84), .B1(n169), .Y(n2469) );
  OA22X1 U2637 ( .A0(n193), .A1(n10960), .B0(n77), .B1(n10950), .Y(n10970) );
  CLKINVX1 U2638 ( .A(stg_reg[136]), .Y(n10960) );
  OA22X1 U2639 ( .A0(n207), .A1(n10900), .B0(n77), .B1(n139), .Y(n10910) );
  CLKINVX1 U2640 ( .A(stg_reg[137]), .Y(n10900) );
  OA22X1 U2641 ( .A0(n199), .A1(n10850), .B0(n75), .B1(n140), .Y(n10860) );
  CLKINVX1 U2642 ( .A(stg_reg[138]), .Y(n10850) );
  OA22X1 U2643 ( .A0(n197), .A1(n10800), .B0(n82), .B1(n145), .Y(n10810) );
  CLKINVX1 U2644 ( .A(stg_reg[139]), .Y(n10800) );
  OA22X1 U2645 ( .A0(n207), .A1(n10750), .B0(n79), .B1(n146), .Y(n10760) );
  CLKINVX1 U2646 ( .A(stg_reg[140]), .Y(n10750) );
  OA22X1 U2647 ( .A0(n199), .A1(n2893), .B0(n77), .B1(n158), .Y(n2399) );
  OA22X1 U2648 ( .A0(n189), .A1(n10700), .B0(n78), .B1(n159), .Y(n10710) );
  CLKINVX1 U2649 ( .A(stg_reg[141]), .Y(n10700) );
  OA22X1 U2650 ( .A0(n195), .A1(n2881), .B0(n84), .B1(n160), .Y(n2395) );
  OA22X1 U2651 ( .A0(n185), .A1(n10650), .B0(n75), .B1(n161), .Y(n10660) );
  CLKINVX1 U2652 ( .A(stg_reg[142]), .Y(n10650) );
  CLKINVX1 U2653 ( .A(stg_reg[145]), .Y(n1271) );
  CLKINVX1 U2654 ( .A(stg_reg[146]), .Y(n1262) );
  CLKINVX1 U2655 ( .A(stg_reg[147]), .Y(n1253) );
  CLKINVX1 U2656 ( .A(stg_reg[148]), .Y(n1244) );
  CLKINVX1 U2657 ( .A(stg_reg[144]), .Y(n1280) );
  AO22X1 U2658 ( .A0(n1575), .A1(n9460), .B0(stg4_img[24]), .B1(n54), .Y(n2267) );
  AO22X1 U2659 ( .A0(n1572), .A1(n9450), .B0(stg4_img[23]), .B1(n62), .Y(n2268) );
  AO22X1 U2660 ( .A0(n1569), .A1(n9410), .B0(stg4_img[22]), .B1(n56), .Y(n2269) );
  AO22X1 U2661 ( .A0(n1566), .A1(n9460), .B0(stg4_img[21]), .B1(n68), .Y(n2270) );
  AO22X1 U2662 ( .A0(n1563), .A1(n9450), .B0(stg4_img[20]), .B1(n58), .Y(n2271) );
  AO22X1 U2663 ( .A0(n1560), .A1(n9410), .B0(stg4_img[19]), .B1(n62), .Y(n2272) );
  AO22X1 U2664 ( .A0(n1557), .A1(n9450), .B0(stg4_img[18]), .B1(n54), .Y(n2273) );
  AO22X1 U2665 ( .A0(n1554), .A1(n9460), .B0(stg4_img[17]), .B1(n68), .Y(n2274) );
  AO22X1 U2666 ( .A0(n1609), .A1(n9440), .B0(stg4_img[8]), .B1(n64), .Y(n2299)
         );
  AO22X1 U2667 ( .A0(n1607), .A1(n9440), .B0(stg4_img[7]), .B1(n72), .Y(n2300)
         );
  AO22X1 U2668 ( .A0(n1605), .A1(n9440), .B0(stg4_img[6]), .B1(n58), .Y(n2301)
         );
  AO22X1 U2669 ( .A0(n1603), .A1(n9450), .B0(stg4_img[5]), .B1(n70), .Y(n2302)
         );
  AO22X1 U2670 ( .A0(n1601), .A1(n9450), .B0(stg4_img[4]), .B1(n54), .Y(n2303)
         );
  AO22X1 U2671 ( .A0(n1599), .A1(n9450), .B0(stg4_img[3]), .B1(n66), .Y(n2304)
         );
  AO22X1 U2672 ( .A0(n1597), .A1(n9450), .B0(stg4_img[2]), .B1(n72), .Y(n2305)
         );
  AO22X1 U2673 ( .A0(n1595), .A1(n9450), .B0(stg4_img[1]), .B1(n72), .Y(n2306)
         );
  AO22X1 U2674 ( .A0(n1470), .A1(n9410), .B0(stg4_img[53]), .B1(n66), .Y(n2206) );
  AO22X1 U2675 ( .A0(n1467), .A1(n9410), .B0(stg4_img[52]), .B1(n60), .Y(n2207) );
  AO22X1 U2676 ( .A0(n1464), .A1(n9420), .B0(stg4_img[51]), .B1(n68), .Y(n2208) );
  AO22X1 U2677 ( .A0(n1461), .A1(n9420), .B0(stg4_img[50]), .B1(n68), .Y(n2209) );
  AO22X1 U2678 ( .A0(n1458), .A1(n9420), .B0(stg4_img[49]), .B1(n56), .Y(n2210) );
  AO22X1 U2679 ( .A0(n1527), .A1(n9430), .B0(stg4_img[40]), .B1(n62), .Y(n2235) );
  AO22X1 U2680 ( .A0(n1524), .A1(n9440), .B0(stg4_img[39]), .B1(n72), .Y(n2236) );
  AO22X1 U2681 ( .A0(n1521), .A1(n9430), .B0(stg4_img[38]), .B1(n60), .Y(n2237) );
  AO22X1 U2682 ( .A0(n1518), .A1(n9440), .B0(stg4_img[37]), .B1(n64), .Y(n2238) );
  AO22X1 U2683 ( .A0(n1515), .A1(n9430), .B0(stg4_img[36]), .B1(n70), .Y(n2239) );
  AO22X1 U2684 ( .A0(n1512), .A1(n9450), .B0(stg4_img[35]), .B1(n62), .Y(n2240) );
  AO22X1 U2685 ( .A0(n1509), .A1(n9410), .B0(stg4_img[34]), .B1(n66), .Y(n2241) );
  AO22X1 U2686 ( .A0(n1506), .A1(n9430), .B0(stg4_img[33]), .B1(n72), .Y(n2242) );
  AO22X1 U2687 ( .A0(n1479), .A1(n9410), .B0(stg4_img[56]), .B1(n66), .Y(n2203) );
  AO22X1 U2688 ( .A0(n1476), .A1(n9410), .B0(stg4_img[55]), .B1(n56), .Y(n2204) );
  AO22X1 U2689 ( .A0(n1473), .A1(n9410), .B0(stg4_img[54]), .B1(n56), .Y(n2205) );
  OA22X1 U2690 ( .A0(n203), .A1(n10600), .B0(n80), .B1(n170), .Y(n10610) );
  CLKINVX1 U2691 ( .A(stg_reg[143]), .Y(n10600) );
  NAND2X1 U2692 ( .A(stg2_real_12__15_), .B(n885), .Y(n2698) );
  CLKINVX1 U2693 ( .A(stg_reg[44]), .Y(n2483) );
  CLKINVX1 U2694 ( .A(stg_reg[45]), .Y(n2478) );
  AND2XL U2695 ( .A(fir_valid), .B(n177), .Y(n10380) );
  CLKINVX1 U2696 ( .A(stg_reg[149]), .Y(n1235) );
  CLKINVX1 U2697 ( .A(stg_reg[150]), .Y(n1226) );
  CLKINVX1 U2698 ( .A(stg_reg[151]), .Y(n1217) );
  CLKINVX1 U2699 ( .A(stg_reg[152]), .Y(n1208) );
  CLKINVX1 U2700 ( .A(stg_reg[153]), .Y(n1199) );
  CLKINVX1 U2701 ( .A(stg_reg[154]), .Y(n1190) );
  CLKINVX1 U2702 ( .A(stg_reg[155]), .Y(n1181) );
  CLKINVX1 U2703 ( .A(stg_reg[59]), .Y(n2595) );
  CLKINVX1 U2704 ( .A(stg_reg[60]), .Y(n2586) );
  CLKINVX1 U2705 ( .A(stg_reg[61]), .Y(n2577) );
  AO22X1 U2706 ( .A0(n1437), .A1(n9420), .B0(stg4_img[48]), .B1(n64), .Y(n2211) );
  AO22X1 U2707 ( .A0(n1581), .A1(n9450), .B0(stg4_img[0]), .B1(n64), .Y(n2307)
         );
  AO22X1 U2708 ( .A0(n1485), .A1(n9430), .B0(stg4_img[32]), .B1(n70), .Y(n2243) );
  AO22X1 U2709 ( .A0(n1533), .A1(n9420), .B0(stg4_img[16]), .B1(n58), .Y(n2275) );
  NAND2X1 U2710 ( .A(stg2_real_12__0_), .B(n880), .Y(n1275) );
  NOR3BXL U2711 ( .AN(fir_valid), .B(n10390), .C(n10480), .Y(N37) );
  AOI21X1 U2712 ( .A0(n9260), .A1(n10410), .B0(n10400), .Y(N38) );
  INVXL U2713 ( .A(fir_valid), .Y(n10400) );
  CLKINVX1 U2714 ( .A(stg_reg[78]), .Y(n3086) );
  CLKINVX1 U2715 ( .A(stg_reg[79]), .Y(n3084) );
  CLKINVX1 U2716 ( .A(stg_reg[46]), .Y(n2473) );
  CLKINVX1 U2717 ( .A(stg_reg[47]), .Y(n2468) );
  CLKINVX1 U2718 ( .A(stg_reg[156]), .Y(n1172) );
  CLKINVX1 U2719 ( .A(stg_reg[157]), .Y(n1163) );
  CLKINVX1 U2720 ( .A(stg_reg[158]), .Y(n1154) );
  CLKINVX1 U2721 ( .A(stg_reg[159]), .Y(n2704) );
  CLKINVX1 U2722 ( .A(stg_reg[62]), .Y(n2568) );
  CLKINVX1 U2723 ( .A(stg_reg[63]), .Y(n2560) );
  CLKINVX1 U2724 ( .A(stg_reg[94]), .Y(n2708) );
  CLKINVX1 U2725 ( .A(stg_reg[95]), .Y(n3068) );
  NAND2X1 U2726 ( .A(n1791), .B(n10190), .Y(n1792) );
  MX2XL U2727 ( .A(fft_d2[0]), .B(n1438), .S0(n10060), .Y(N919) );
  MX2XL U2728 ( .A(fft_d6[0]), .B(n1534), .S0(n9980), .Y(N983) );
  MX2XL U2729 ( .A(fft_d10[0]), .B(n1486), .S0(n9910), .Y(N951) );
  MX2XL U2730 ( .A(fft_d14[0]), .B(n1582), .S0(n9840), .Y(N1015) );
  MX2XL U2731 ( .A(fft_d2[1]), .B(n1459), .S0(n10060), .Y(N920) );
  MX2XL U2732 ( .A(fft_d6[1]), .B(n1555), .S0(n9980), .Y(N984) );
  MX2XL U2733 ( .A(fft_d10[1]), .B(n1507), .S0(n9910), .Y(N952) );
  MX2XL U2734 ( .A(fft_d14[1]), .B(n1596), .S0(n9840), .Y(N1016) );
  MX2XL U2735 ( .A(fft_d2[2]), .B(n1462), .S0(n10060), .Y(N921) );
  MX2XL U2736 ( .A(fft_d6[2]), .B(n1558), .S0(n9980), .Y(N985) );
  MX2XL U2737 ( .A(fft_d10[2]), .B(n1510), .S0(n9910), .Y(N953) );
  MX2XL U2738 ( .A(fft_d14[2]), .B(n1598), .S0(n9840), .Y(N1017) );
  MX2XL U2739 ( .A(fft_d2[3]), .B(n1465), .S0(n10060), .Y(N922) );
  MX2XL U2740 ( .A(fft_d6[3]), .B(n1561), .S0(n9990), .Y(N986) );
  MX2XL U2741 ( .A(fft_d10[3]), .B(n1513), .S0(n9910), .Y(N954) );
  MX2XL U2742 ( .A(fft_d14[3]), .B(n1600), .S0(n9840), .Y(N1018) );
  MX2XL U2743 ( .A(fft_d2[4]), .B(n1468), .S0(n10060), .Y(N923) );
  MX2XL U2744 ( .A(fft_d6[4]), .B(n1564), .S0(n9990), .Y(N987) );
  MX2XL U2745 ( .A(fft_d10[4]), .B(n1516), .S0(n9910), .Y(N955) );
  MX2XL U2746 ( .A(fft_d14[4]), .B(n1602), .S0(n9840), .Y(N1019) );
  MX2XL U2747 ( .A(fft_d2[5]), .B(n1471), .S0(n10060), .Y(N924) );
  MX2XL U2748 ( .A(fft_d6[5]), .B(n1567), .S0(n9990), .Y(N988) );
  MX2XL U2749 ( .A(fft_d10[5]), .B(n1519), .S0(n9910), .Y(N956) );
  MX2XL U2750 ( .A(fft_d14[5]), .B(n1604), .S0(n9840), .Y(N1020) );
  MX2XL U2751 ( .A(fft_d2[6]), .B(n1474), .S0(n10060), .Y(N925) );
  MX2XL U2752 ( .A(fft_d6[6]), .B(n1570), .S0(n9990), .Y(N989) );
  MX2XL U2753 ( .A(fft_d10[6]), .B(n1522), .S0(n9910), .Y(N957) );
  MX2XL U2754 ( .A(fft_d14[6]), .B(n1606), .S0(n9840), .Y(N1021) );
  MX2XL U2755 ( .A(fft_d2[7]), .B(n1477), .S0(n10060), .Y(N926) );
  MX2XL U2756 ( .A(fft_d6[7]), .B(n1573), .S0(n9990), .Y(N990) );
  MX2XL U2757 ( .A(fft_d10[7]), .B(n1525), .S0(n9910), .Y(N958) );
  MX2XL U2758 ( .A(fft_d14[7]), .B(n1608), .S0(n9840), .Y(N1022) );
  MX2XL U2759 ( .A(fft_d2[8]), .B(n1480), .S0(n10060), .Y(N927) );
  MX2XL U2760 ( .A(fft_d6[8]), .B(n1576), .S0(n9990), .Y(N991) );
  MX2XL U2761 ( .A(fft_d10[8]), .B(n1528), .S0(n9920), .Y(N959) );
  MX2XL U2762 ( .A(fft_d14[8]), .B(n1610), .S0(n9840), .Y(N1023) );
  MX2XL U2763 ( .A(fft_d2[9]), .B(n1483), .S0(n10060), .Y(N928) );
  MX2XL U2764 ( .A(fft_d6[9]), .B(n1579), .S0(n9990), .Y(N992) );
  MX2XL U2765 ( .A(fft_d10[9]), .B(n1531), .S0(n9920), .Y(N960) );
  MX2XL U2766 ( .A(fft_d14[9]), .B(n1612), .S0(n9840), .Y(N1024) );
  MX2XL U2767 ( .A(fft_d2[10]), .B(n1441), .S0(n10060), .Y(N929) );
  MX2XL U2768 ( .A(fft_d6[10]), .B(n1537), .S0(n9990), .Y(N993) );
  MX2XL U2769 ( .A(fft_d10[10]), .B(n1489), .S0(n9920), .Y(N961) );
  MX2XL U2770 ( .A(fft_d14[10]), .B(n1584), .S0(n9840), .Y(N1025) );
  MX2XL U2771 ( .A(fft_d2[11]), .B(n1444), .S0(n10070), .Y(N930) );
  MX2XL U2772 ( .A(fft_d6[11]), .B(n1540), .S0(n9990), .Y(N994) );
  MX2XL U2773 ( .A(fft_d10[11]), .B(n1492), .S0(n9920), .Y(N962) );
  MX2XL U2774 ( .A(fft_d14[11]), .B(n1586), .S0(n9840), .Y(N1026) );
  MX2XL U2775 ( .A(fft_d2[12]), .B(n1447), .S0(n10070), .Y(N931) );
  MX2XL U2776 ( .A(fft_d6[12]), .B(n1543), .S0(n9990), .Y(N995) );
  MX2XL U2777 ( .A(fft_d10[12]), .B(n1495), .S0(n9920), .Y(N963) );
  MX2XL U2778 ( .A(fft_d14[12]), .B(n1588), .S0(n9840), .Y(N1027) );
  MX2XL U2779 ( .A(fft_d2[13]), .B(n1450), .S0(n10070), .Y(N932) );
  MX2XL U2780 ( .A(fft_d6[13]), .B(n1546), .S0(n9990), .Y(N996) );
  MX2XL U2781 ( .A(fft_d10[13]), .B(n1498), .S0(n9920), .Y(N964) );
  MX2XL U2782 ( .A(fft_d14[13]), .B(n1590), .S0(n9850), .Y(N1028) );
  MX2XL U2783 ( .A(fft_d2[14]), .B(n1453), .S0(n10070), .Y(N933) );
  MX2XL U2784 ( .A(fft_d6[14]), .B(n1549), .S0(n9990), .Y(N997) );
  MX2XL U2785 ( .A(fft_d10[14]), .B(n1501), .S0(n9920), .Y(N965) );
  MX2XL U2786 ( .A(fft_d14[14]), .B(n1592), .S0(n9850), .Y(N1029) );
  MX2XL U2787 ( .A(fft_d2[15]), .B(n1456), .S0(n10070), .Y(N934) );
  MX2XL U2788 ( .A(fft_d6[15]), .B(n1552), .S0(n9990), .Y(N998) );
  MX2XL U2789 ( .A(fft_d10[15]), .B(n1504), .S0(n9920), .Y(N966) );
  MX2XL U2790 ( .A(fft_d14[15]), .B(n1594), .S0(n9850), .Y(N1030) );
  MX2XL U2791 ( .A(fft_d2[16]), .B(n1614), .S0(n10070), .Y(N935) );
  MX2XL U2792 ( .A(fft_d6[16]), .B(n1710), .S0(n10000), .Y(N999) );
  MX2XL U2793 ( .A(fft_d10[16]), .B(n1662), .S0(n9920), .Y(N967) );
  MX2XL U2794 ( .A(fft_d14[16]), .B(n1758), .S0(n9850), .Y(N1031) );
  MX2XL U2795 ( .A(fft_d2[17]), .B(n1635), .S0(n10070), .Y(N936) );
  MX2XL U2796 ( .A(fft_d6[17]), .B(n1731), .S0(n10000), .Y(N1000) );
  MX2XL U2797 ( .A(fft_d10[17]), .B(n1683), .S0(n9920), .Y(N968) );
  MX2XL U2798 ( .A(fft_d14[17]), .B(n1772), .S0(n9850), .Y(N1032) );
  MX2XL U2799 ( .A(fft_d2[18]), .B(n1638), .S0(n10070), .Y(N937) );
  MX2XL U2800 ( .A(fft_d6[18]), .B(n1734), .S0(n10000), .Y(N1001) );
  MX2XL U2801 ( .A(fft_d10[18]), .B(n1686), .S0(n9920), .Y(N969) );
  MX2XL U2802 ( .A(fft_d14[18]), .B(n1774), .S0(n9850), .Y(N1033) );
  MX2XL U2803 ( .A(fft_d2[19]), .B(n1641), .S0(n10070), .Y(N938) );
  MX2XL U2804 ( .A(fft_d6[19]), .B(n1737), .S0(n10000), .Y(N1002) );
  MX2XL U2805 ( .A(fft_d10[19]), .B(n1689), .S0(n9920), .Y(N970) );
  MX2XL U2806 ( .A(fft_d14[19]), .B(n1776), .S0(n9850), .Y(N1034) );
  MX2XL U2807 ( .A(fft_d2[20]), .B(n1644), .S0(n10070), .Y(N939) );
  MX2XL U2808 ( .A(fft_d6[20]), .B(n1740), .S0(n10000), .Y(N1003) );
  MX2XL U2809 ( .A(fft_d10[20]), .B(n1692), .S0(n9920), .Y(N971) );
  MX2XL U2810 ( .A(fft_d14[20]), .B(n1778), .S0(n9850), .Y(N1035) );
  MX2XL U2811 ( .A(fft_d2[21]), .B(n1647), .S0(n10070), .Y(N940) );
  MX2XL U2812 ( .A(fft_d6[21]), .B(n1743), .S0(n10000), .Y(N1004) );
  MX2XL U2813 ( .A(fft_d10[21]), .B(n1695), .S0(n9930), .Y(N972) );
  MX2XL U2814 ( .A(fft_d14[21]), .B(n1780), .S0(n9850), .Y(N1036) );
  MX2XL U2815 ( .A(fft_d2[22]), .B(n1650), .S0(n10070), .Y(N941) );
  MX2XL U2816 ( .A(fft_d6[22]), .B(n1746), .S0(n10000), .Y(N1005) );
  MX2XL U2817 ( .A(fft_d10[22]), .B(n1698), .S0(n9930), .Y(N973) );
  MX2XL U2818 ( .A(fft_d14[22]), .B(n1782), .S0(n9850), .Y(N1037) );
  MX2XL U2819 ( .A(fft_d2[23]), .B(n1653), .S0(n10070), .Y(N942) );
  MX2XL U2820 ( .A(fft_d6[23]), .B(n1749), .S0(n10000), .Y(N1006) );
  MX2XL U2821 ( .A(fft_d10[23]), .B(n1701), .S0(n9930), .Y(N974) );
  MX2XL U2822 ( .A(fft_d14[23]), .B(n1784), .S0(n9850), .Y(N1038) );
  MX2XL U2823 ( .A(fft_d2[24]), .B(n1656), .S0(n10080), .Y(N943) );
  MX2XL U2824 ( .A(fft_d6[24]), .B(n1752), .S0(n10000), .Y(N1007) );
  MX2XL U2825 ( .A(fft_d10[24]), .B(n1704), .S0(n9930), .Y(N975) );
  MX2XL U2826 ( .A(fft_d14[24]), .B(n1786), .S0(n9850), .Y(N1039) );
  MX2XL U2827 ( .A(fft_d2[25]), .B(n1659), .S0(n10080), .Y(N944) );
  MX2XL U2828 ( .A(fft_d6[25]), .B(n1755), .S0(n10000), .Y(N1008) );
  MX2XL U2829 ( .A(fft_d10[25]), .B(n1707), .S0(n9930), .Y(N976) );
  MX2XL U2830 ( .A(fft_d14[25]), .B(n1788), .S0(n9850), .Y(N1040) );
  MX2XL U2831 ( .A(fft_d2[26]), .B(n1617), .S0(n10080), .Y(N945) );
  MX2XL U2832 ( .A(fft_d6[26]), .B(n1713), .S0(n10000), .Y(N1009) );
  MX2XL U2833 ( .A(fft_d10[26]), .B(n1665), .S0(n9930), .Y(N977) );
  MX2XL U2834 ( .A(fft_d14[26]), .B(n1760), .S0(n9860), .Y(N1041) );
  MX2XL U2835 ( .A(fft_d2[27]), .B(n1620), .S0(n10080), .Y(N946) );
  MX2XL U2836 ( .A(fft_d6[27]), .B(n1716), .S0(n10000), .Y(N1010) );
  MX2XL U2837 ( .A(fft_d10[27]), .B(n1668), .S0(n9930), .Y(N978) );
  MX2XL U2838 ( .A(fft_d14[27]), .B(n1762), .S0(n9860), .Y(N1042) );
  MX2XL U2839 ( .A(fft_d2[28]), .B(n1623), .S0(n10080), .Y(N947) );
  MX2XL U2840 ( .A(fft_d6[28]), .B(n1719), .S0(n10000), .Y(N1011) );
  MX2XL U2841 ( .A(fft_d10[28]), .B(n1671), .S0(n9930), .Y(N979) );
  MX2XL U2842 ( .A(fft_d14[28]), .B(n1764), .S0(n9860), .Y(N1043) );
  MX2XL U2843 ( .A(fft_d2[29]), .B(n1626), .S0(n10080), .Y(N948) );
  MX2XL U2844 ( .A(fft_d6[29]), .B(n1722), .S0(n10010), .Y(N1012) );
  MX2XL U2845 ( .A(fft_d10[29]), .B(n1674), .S0(n9930), .Y(N980) );
  MX2XL U2846 ( .A(fft_d14[29]), .B(n1766), .S0(n9860), .Y(N1044) );
  MX2XL U2847 ( .A(fft_d2[30]), .B(n1629), .S0(n10080), .Y(N949) );
  MX2XL U2848 ( .A(fft_d6[30]), .B(n1725), .S0(n10010), .Y(N1013) );
  MX2XL U2849 ( .A(fft_d10[30]), .B(n1677), .S0(n9930), .Y(N981) );
  MX2XL U2850 ( .A(fft_d14[30]), .B(n1768), .S0(n9860), .Y(N1045) );
  MX2XL U2851 ( .A(fft_d2[31]), .B(n1632), .S0(n10080), .Y(N950) );
  MX2XL U2852 ( .A(fft_d6[31]), .B(n1728), .S0(n10010), .Y(N1014) );
  MX2XL U2853 ( .A(fft_d10[31]), .B(n1680), .S0(n9930), .Y(N982) );
  MX2XL U2854 ( .A(fft_d14[31]), .B(n1770), .S0(n9860), .Y(N1046) );
  MX2XL U2855 ( .A(fft_d1[16]), .B(n1613), .S0(n10090), .Y(N679) );
  MX2XL U2856 ( .A(fft_d1[0]), .B(n1437), .S0(n10080), .Y(N663) );
  MX2XL U2857 ( .A(fft_d1[2]), .B(n1461), .S0(n10080), .Y(N665) );
  MX2XL U2858 ( .A(fft_d1[18]), .B(n1637), .S0(n10100), .Y(N681) );
  MX2XL U2859 ( .A(fft_d4[0]), .B(n1439), .S0(n10030), .Y(N1047) );
  MX2XL U2860 ( .A(fft_d5[0]), .B(n1533), .S0(n10010), .Y(N727) );
  MX2XL U2861 ( .A(fft_d8[0]), .B(n1535), .S0(n9960), .Y(N1111) );
  MX2XL U2862 ( .A(fft_d9[0]), .B(n1485), .S0(n9930), .Y(N695) );
  MX2XL U2863 ( .A(fft_d12[0]), .B(n1487), .S0(n9880), .Y(N1079) );
  MX2XL U2864 ( .A(fft_d13[0]), .B(n1581), .S0(n9860), .Y(N759) );
  MX2XL U2865 ( .A(fft_d1[1]), .B(n1458), .S0(n10080), .Y(N664) );
  MX2XL U2866 ( .A(fft_d4[1]), .B(n1460), .S0(n10030), .Y(N1048) );
  MX2XL U2867 ( .A(fft_d5[1]), .B(n1554), .S0(n10010), .Y(N728) );
  MX2XL U2868 ( .A(fft_d8[1]), .B(n1556), .S0(n9960), .Y(N1112) );
  MX2XL U2869 ( .A(fft_d9[1]), .B(n1506), .S0(n9930), .Y(N696) );
  MX2XL U2870 ( .A(fft_d12[1]), .B(n1508), .S0(n9890), .Y(N1080) );
  MX2XL U2871 ( .A(fft_d13[1]), .B(n1595), .S0(n9860), .Y(N760) );
  MX2XL U2872 ( .A(fft_d4[2]), .B(n1463), .S0(n10030), .Y(N1049) );
  MX2XL U2873 ( .A(fft_d5[2]), .B(n1557), .S0(n10010), .Y(N729) );
  MX2XL U2874 ( .A(fft_d8[2]), .B(n1559), .S0(n9960), .Y(N1113) );
  MX2XL U2875 ( .A(fft_d9[2]), .B(n1509), .S0(n9940), .Y(N697) );
  MX2XL U2876 ( .A(fft_d12[2]), .B(n1511), .S0(n9890), .Y(N1081) );
  MX2XL U2877 ( .A(fft_d13[2]), .B(n1597), .S0(n9860), .Y(N761) );
  MX2XL U2878 ( .A(fft_d1[3]), .B(n1464), .S0(n10080), .Y(N666) );
  MX2XL U2879 ( .A(fft_d4[3]), .B(n1466), .S0(n10030), .Y(N1050) );
  MX2XL U2880 ( .A(fft_d5[3]), .B(n1560), .S0(n10010), .Y(N730) );
  MX2XL U2881 ( .A(fft_d8[3]), .B(n1562), .S0(n9960), .Y(N1114) );
  MX2XL U2882 ( .A(fft_d9[3]), .B(n1512), .S0(n9940), .Y(N698) );
  MX2XL U2883 ( .A(fft_d12[3]), .B(n1514), .S0(n9890), .Y(N1082) );
  MX2XL U2884 ( .A(fft_d13[3]), .B(n1599), .S0(n9860), .Y(N762) );
  MX2XL U2885 ( .A(fft_d1[4]), .B(n1467), .S0(n10080), .Y(N667) );
  MX2XL U2886 ( .A(fft_d4[4]), .B(n1469), .S0(n10040), .Y(N1051) );
  MX2XL U2887 ( .A(fft_d5[4]), .B(n1563), .S0(n10010), .Y(N731) );
  MX2XL U2888 ( .A(fft_d8[4]), .B(n1565), .S0(n9960), .Y(N1115) );
  MX2XL U2889 ( .A(fft_d9[4]), .B(n1515), .S0(n9940), .Y(N699) );
  MX2XL U2890 ( .A(fft_d12[4]), .B(n1517), .S0(n9890), .Y(N1083) );
  MX2XL U2891 ( .A(fft_d13[4]), .B(n1601), .S0(n9860), .Y(N763) );
  MX2XL U2892 ( .A(fft_d1[5]), .B(n1470), .S0(n10090), .Y(N668) );
  MX2XL U2893 ( .A(fft_d4[5]), .B(n1472), .S0(n10040), .Y(N1052) );
  MX2XL U2894 ( .A(fft_d5[5]), .B(n1566), .S0(n10010), .Y(N732) );
  MX2XL U2895 ( .A(fft_d8[5]), .B(n1568), .S0(n9960), .Y(N1116) );
  MX2XL U2896 ( .A(fft_d9[5]), .B(n1518), .S0(n9940), .Y(N700) );
  MX2XL U2897 ( .A(fft_d12[5]), .B(n1520), .S0(n9890), .Y(N1084) );
  MX2XL U2898 ( .A(fft_d13[5]), .B(n1603), .S0(n9860), .Y(N764) );
  MX2XL U2899 ( .A(fft_d1[6]), .B(n1473), .S0(n10090), .Y(N669) );
  MX2XL U2900 ( .A(fft_d4[6]), .B(n1475), .S0(n10040), .Y(N1053) );
  MX2XL U2901 ( .A(fft_d5[6]), .B(n1569), .S0(n10010), .Y(N733) );
  MX2XL U2902 ( .A(fft_d8[6]), .B(n1571), .S0(n9960), .Y(N1117) );
  MX2XL U2903 ( .A(fft_d9[6]), .B(n1521), .S0(n9940), .Y(N701) );
  MX2XL U2904 ( .A(fft_d12[6]), .B(n1523), .S0(n9890), .Y(N1085) );
  MX2XL U2905 ( .A(fft_d13[6]), .B(n1605), .S0(n9860), .Y(N765) );
  MX2XL U2906 ( .A(fft_d1[7]), .B(n1476), .S0(n10090), .Y(N670) );
  MX2XL U2907 ( .A(fft_d4[7]), .B(n1478), .S0(n10040), .Y(N1054) );
  MX2XL U2908 ( .A(fft_d5[7]), .B(n1572), .S0(n10010), .Y(N734) );
  MX2XL U2909 ( .A(fft_d8[7]), .B(n1574), .S0(n9960), .Y(N1118) );
  MX2XL U2910 ( .A(fft_d9[7]), .B(n1524), .S0(n9940), .Y(N702) );
  MX2XL U2911 ( .A(fft_d12[7]), .B(n1526), .S0(n9890), .Y(N1086) );
  MX2XL U2912 ( .A(fft_d13[7]), .B(n1607), .S0(n9870), .Y(N766) );
  MX2XL U2913 ( .A(fft_d1[8]), .B(n1479), .S0(n10090), .Y(N671) );
  MX2XL U2914 ( .A(fft_d4[8]), .B(n1481), .S0(n10040), .Y(N1055) );
  MX2XL U2915 ( .A(fft_d5[8]), .B(n1575), .S0(n10010), .Y(N735) );
  MX2XL U2916 ( .A(fft_d8[8]), .B(n1577), .S0(n9960), .Y(N1119) );
  MX2XL U2917 ( .A(fft_d9[8]), .B(n1527), .S0(n9940), .Y(N703) );
  MX2XL U2918 ( .A(fft_d12[8]), .B(n1529), .S0(n9890), .Y(N1087) );
  MX2XL U2919 ( .A(fft_d13[8]), .B(n1609), .S0(n9870), .Y(N767) );
  MX2XL U2920 ( .A(fft_d1[9]), .B(n1482), .S0(n10090), .Y(N672) );
  MX2XL U2921 ( .A(fft_d4[9]), .B(n1484), .S0(n10040), .Y(N1056) );
  MX2XL U2922 ( .A(fft_d5[9]), .B(n1578), .S0(n10010), .Y(N736) );
  MX2XL U2923 ( .A(fft_d8[9]), .B(n1580), .S0(n9970), .Y(N1120) );
  MX2XL U2924 ( .A(fft_d9[9]), .B(n1530), .S0(n9940), .Y(N704) );
  MX2XL U2925 ( .A(fft_d12[9]), .B(n1532), .S0(n9890), .Y(N1088) );
  MX2XL U2926 ( .A(fft_d13[9]), .B(n1611), .S0(n9870), .Y(N768) );
  MX2XL U2927 ( .A(fft_d1[10]), .B(n1440), .S0(n10090), .Y(N673) );
  MX2XL U2928 ( .A(fft_d4[10]), .B(n1442), .S0(n10040), .Y(N1057) );
  MX2XL U2929 ( .A(fft_d5[10]), .B(n1536), .S0(n10020), .Y(N737) );
  MX2XL U2930 ( .A(fft_d8[10]), .B(n1538), .S0(n9970), .Y(N1121) );
  MX2XL U2931 ( .A(fft_d9[10]), .B(n1488), .S0(n9940), .Y(N705) );
  MX2XL U2932 ( .A(fft_d12[10]), .B(n1490), .S0(n9890), .Y(N1089) );
  MX2XL U2933 ( .A(fft_d13[10]), .B(n1583), .S0(n9870), .Y(N769) );
  MX2XL U2934 ( .A(fft_d1[11]), .B(n1443), .S0(n10090), .Y(N674) );
  MX2XL U2935 ( .A(fft_d4[11]), .B(n1445), .S0(n10040), .Y(N1058) );
  MX2XL U2936 ( .A(fft_d5[11]), .B(n1539), .S0(n10020), .Y(N738) );
  MX2XL U2937 ( .A(fft_d8[11]), .B(n1541), .S0(n9970), .Y(N1122) );
  MX2XL U2938 ( .A(fft_d9[11]), .B(n1491), .S0(n9940), .Y(N706) );
  MX2XL U2939 ( .A(fft_d12[11]), .B(n1493), .S0(n9890), .Y(N1090) );
  MX2XL U2940 ( .A(fft_d13[11]), .B(n1585), .S0(n9870), .Y(N770) );
  MX2XL U2941 ( .A(fft_d1[12]), .B(n1446), .S0(n10090), .Y(N675) );
  MX2XL U2942 ( .A(fft_d4[12]), .B(n1448), .S0(n10040), .Y(N1059) );
  MX2XL U2943 ( .A(fft_d5[12]), .B(n1542), .S0(n10020), .Y(N739) );
  MX2XL U2944 ( .A(fft_d8[12]), .B(n1544), .S0(n9970), .Y(N1123) );
  MX2XL U2945 ( .A(fft_d9[12]), .B(n1494), .S0(n9940), .Y(N707) );
  MX2XL U2946 ( .A(fft_d12[12]), .B(n1496), .S0(n9890), .Y(N1091) );
  MX2XL U2947 ( .A(fft_d13[12]), .B(n1587), .S0(n9870), .Y(N771) );
  MX2XL U2948 ( .A(fft_d1[13]), .B(n1449), .S0(n10090), .Y(N676) );
  MX2XL U2949 ( .A(fft_d4[13]), .B(n1451), .S0(n10040), .Y(N1060) );
  MX2XL U2950 ( .A(fft_d5[13]), .B(n1545), .S0(n10020), .Y(N740) );
  MX2XL U2951 ( .A(fft_d8[13]), .B(n1547), .S0(n9970), .Y(N1124) );
  MX2XL U2952 ( .A(fft_d9[13]), .B(n1497), .S0(n9940), .Y(N708) );
  MX2XL U2953 ( .A(fft_d12[13]), .B(n1499), .S0(n9890), .Y(N1092) );
  MX2XL U2954 ( .A(fft_d13[13]), .B(n1589), .S0(n9870), .Y(N772) );
  MX2XL U2955 ( .A(fft_d1[14]), .B(n1452), .S0(n10090), .Y(N677) );
  MX2XL U2956 ( .A(fft_d4[14]), .B(n1454), .S0(n10040), .Y(N1061) );
  MX2XL U2957 ( .A(fft_d5[14]), .B(n1548), .S0(n10020), .Y(N741) );
  MX2XL U2958 ( .A(fft_d8[14]), .B(n1550), .S0(n9970), .Y(N1125) );
  MX2XL U2959 ( .A(fft_d9[14]), .B(n1500), .S0(n9940), .Y(N709) );
  MX2XL U2960 ( .A(fft_d12[14]), .B(n1502), .S0(n9900), .Y(N1093) );
  MX2XL U2961 ( .A(fft_d13[14]), .B(n1591), .S0(n9870), .Y(N773) );
  MX2XL U2962 ( .A(fft_d1[15]), .B(n1455), .S0(n10090), .Y(N678) );
  MX2XL U2963 ( .A(fft_d4[15]), .B(n1457), .S0(n10040), .Y(N1062) );
  MX2XL U2964 ( .A(fft_d5[15]), .B(n1551), .S0(n10020), .Y(N742) );
  MX2XL U2965 ( .A(fft_d8[15]), .B(n1553), .S0(n9970), .Y(N1126) );
  MX2XL U2966 ( .A(fft_d9[15]), .B(n1503), .S0(n9950), .Y(N710) );
  MX2XL U2967 ( .A(fft_d12[15]), .B(n1505), .S0(n9900), .Y(N1094) );
  MX2XL U2968 ( .A(fft_d13[15]), .B(n1593), .S0(n9870), .Y(N774) );
  MX2XL U2969 ( .A(fft_d4[16]), .B(n1615), .S0(n10040), .Y(N1063) );
  MX2XL U2970 ( .A(fft_d5[16]), .B(n1709), .S0(n10020), .Y(N743) );
  MX2XL U2971 ( .A(fft_d8[16]), .B(n1711), .S0(n9970), .Y(N1127) );
  MX2XL U2972 ( .A(fft_d9[16]), .B(n1661), .S0(n9950), .Y(N711) );
  MX2XL U2973 ( .A(fft_d12[16]), .B(n1663), .S0(n9900), .Y(N1095) );
  MX2XL U2974 ( .A(fft_d13[16]), .B(n1757), .S0(n9870), .Y(N775) );
  MX2XL U2975 ( .A(fft_d1[17]), .B(n1634), .S0(n10090), .Y(N680) );
  MX2XL U2976 ( .A(fft_d4[17]), .B(n1636), .S0(n10050), .Y(N1064) );
  MX2XL U2977 ( .A(fft_d5[17]), .B(n1730), .S0(n10020), .Y(N744) );
  MX2XL U2978 ( .A(fft_d8[17]), .B(n1732), .S0(n9970), .Y(N1128) );
  MX2XL U2979 ( .A(fft_d9[17]), .B(n1682), .S0(n9950), .Y(N712) );
  MX2XL U2980 ( .A(fft_d12[17]), .B(n1684), .S0(n9900), .Y(N1096) );
  MX2XL U2981 ( .A(fft_d13[17]), .B(n1771), .S0(n9870), .Y(N776) );
  MX2XL U2982 ( .A(fft_d4[18]), .B(n1639), .S0(n10050), .Y(N1065) );
  MX2XL U2983 ( .A(fft_d5[18]), .B(n1733), .S0(n10020), .Y(N745) );
  MX2XL U2984 ( .A(fft_d8[18]), .B(n1735), .S0(n9970), .Y(N1129) );
  MX2XL U2985 ( .A(fft_d9[18]), .B(n1685), .S0(n9950), .Y(N713) );
  MX2XL U2986 ( .A(fft_d12[18]), .B(n1687), .S0(n9900), .Y(N1097) );
  MX2XL U2987 ( .A(fft_d13[18]), .B(n1773), .S0(n9870), .Y(N777) );
  MX2XL U2988 ( .A(fft_d1[19]), .B(n1640), .S0(n10100), .Y(N682) );
  MX2XL U2989 ( .A(fft_d4[19]), .B(n1642), .S0(n10050), .Y(N1066) );
  MX2XL U2990 ( .A(fft_d5[19]), .B(n1736), .S0(n10020), .Y(N746) );
  MX2XL U2991 ( .A(fft_d8[19]), .B(n1738), .S0(n9970), .Y(N1130) );
  MX2XL U2992 ( .A(fft_d9[19]), .B(n1688), .S0(n9950), .Y(N714) );
  MX2XL U2993 ( .A(fft_d12[19]), .B(n1690), .S0(n9900), .Y(N1098) );
  MX2XL U2994 ( .A(fft_d13[19]), .B(n1775), .S0(n9870), .Y(N778) );
  MX2XL U2995 ( .A(fft_d1[20]), .B(n1643), .S0(n10100), .Y(N683) );
  MX2XL U2996 ( .A(fft_d4[20]), .B(n1645), .S0(n10050), .Y(N1067) );
  MX2XL U2997 ( .A(fft_d5[20]), .B(n1739), .S0(n10020), .Y(N747) );
  MX2XL U2998 ( .A(fft_d8[20]), .B(n1741), .S0(n9970), .Y(N1131) );
  MX2XL U2999 ( .A(fft_d9[20]), .B(n1691), .S0(n9950), .Y(N715) );
  MX2XL U3000 ( .A(fft_d12[20]), .B(n1693), .S0(n9900), .Y(N1099) );
  MX2XL U3001 ( .A(fft_d13[20]), .B(n1777), .S0(n9880), .Y(N779) );
  MX2XL U3002 ( .A(fft_d1[21]), .B(n1646), .S0(n10100), .Y(N684) );
  MX2XL U3003 ( .A(fft_d4[21]), .B(n1648), .S0(n10050), .Y(N1068) );
  MX2XL U3004 ( .A(fft_d5[21]), .B(n1742), .S0(n10020), .Y(N748) );
  MX2XL U3005 ( .A(fft_d8[21]), .B(n1744), .S0(n9970), .Y(N1132) );
  MX2XL U3006 ( .A(fft_d9[21]), .B(n1694), .S0(n9950), .Y(N716) );
  MX2XL U3007 ( .A(fft_d12[21]), .B(n1696), .S0(n9900), .Y(N1100) );
  MX2XL U3008 ( .A(fft_d13[21]), .B(n1779), .S0(n9880), .Y(N780) );
  MX2XL U3009 ( .A(fft_d1[22]), .B(n1649), .S0(n10100), .Y(N685) );
  MX2XL U3010 ( .A(fft_d4[22]), .B(n1651), .S0(n10050), .Y(N1069) );
  MX2XL U3011 ( .A(fft_d5[22]), .B(n1745), .S0(n10020), .Y(N749) );
  MX2XL U3012 ( .A(fft_d8[22]), .B(n1747), .S0(n9980), .Y(N1133) );
  MX2XL U3013 ( .A(fft_d9[22]), .B(n1697), .S0(n9950), .Y(N717) );
  MX2XL U3014 ( .A(fft_d12[22]), .B(n1699), .S0(n9900), .Y(N1101) );
  MX2XL U3015 ( .A(fft_d13[22]), .B(n1781), .S0(n9880), .Y(N781) );
  MX2XL U3016 ( .A(fft_d1[23]), .B(n1652), .S0(n10100), .Y(N686) );
  MX2XL U3017 ( .A(fft_d4[23]), .B(n1654), .S0(n10050), .Y(N1070) );
  MX2XL U3018 ( .A(fft_d5[23]), .B(n1748), .S0(n10030), .Y(N750) );
  MX2XL U3019 ( .A(fft_d8[23]), .B(n1750), .S0(n9980), .Y(N1134) );
  MX2XL U3020 ( .A(fft_d9[23]), .B(n1700), .S0(n9950), .Y(N718) );
  MX2XL U3021 ( .A(fft_d12[23]), .B(n1702), .S0(n9900), .Y(N1102) );
  MX2XL U3022 ( .A(fft_d13[23]), .B(n1783), .S0(n9880), .Y(N782) );
  MX2XL U3023 ( .A(fft_d1[24]), .B(n1655), .S0(n10100), .Y(N687) );
  MX2XL U3024 ( .A(fft_d4[24]), .B(n1657), .S0(n10050), .Y(N1071) );
  MX2XL U3025 ( .A(fft_d5[24]), .B(n1751), .S0(n10030), .Y(N751) );
  MX2XL U3026 ( .A(fft_d8[24]), .B(n1753), .S0(n9980), .Y(N1135) );
  MX2XL U3027 ( .A(fft_d9[24]), .B(n1703), .S0(n9950), .Y(N719) );
  MX2XL U3028 ( .A(fft_d12[24]), .B(n1705), .S0(n9900), .Y(N1103) );
  MX2XL U3029 ( .A(fft_d13[24]), .B(n1785), .S0(n9880), .Y(N783) );
  MX2XL U3030 ( .A(fft_d1[25]), .B(n1658), .S0(n10100), .Y(N688) );
  MX2XL U3031 ( .A(fft_d4[25]), .B(n1660), .S0(n10050), .Y(N1072) );
  MX2XL U3032 ( .A(fft_d5[25]), .B(n1754), .S0(n10030), .Y(N752) );
  MX2XL U3033 ( .A(fft_d8[25]), .B(n1756), .S0(n9980), .Y(N1136) );
  MX2XL U3034 ( .A(fft_d9[25]), .B(n1706), .S0(n9950), .Y(N720) );
  MX2XL U3035 ( .A(fft_d12[25]), .B(n1708), .S0(n9900), .Y(N1104) );
  MX2XL U3036 ( .A(fft_d13[25]), .B(n1787), .S0(n9880), .Y(N784) );
  MX2XL U3037 ( .A(fft_d1[26]), .B(n1616), .S0(n10100), .Y(N689) );
  MX2XL U3038 ( .A(fft_d4[26]), .B(n1618), .S0(n10050), .Y(N1073) );
  MX2XL U3039 ( .A(fft_d5[26]), .B(n1712), .S0(n10030), .Y(N753) );
  MX2XL U3040 ( .A(fft_d8[26]), .B(n1714), .S0(n9980), .Y(N1137) );
  MX2XL U3041 ( .A(fft_d9[26]), .B(n1664), .S0(n9950), .Y(N721) );
  MX2XL U3042 ( .A(fft_d12[26]), .B(n1666), .S0(n9900), .Y(N1105) );
  MX2XL U3043 ( .A(fft_d13[26]), .B(n1759), .S0(n9880), .Y(N785) );
  MX2XL U3044 ( .A(fft_d1[27]), .B(n1619), .S0(n10100), .Y(N690) );
  MX2XL U3045 ( .A(fft_d4[27]), .B(n1621), .S0(n10050), .Y(N1074) );
  MX2XL U3046 ( .A(fft_d5[27]), .B(n1715), .S0(n10030), .Y(N754) );
  MX2XL U3047 ( .A(fft_d8[27]), .B(n1717), .S0(n9980), .Y(N1138) );
  MX2XL U3048 ( .A(fft_d9[27]), .B(n1667), .S0(n9950), .Y(N722) );
  MX2XL U3049 ( .A(fft_d12[27]), .B(n1669), .S0(n9910), .Y(N1106) );
  MX2XL U3050 ( .A(fft_d13[27]), .B(n1761), .S0(n9880), .Y(N786) );
  MX2XL U3051 ( .A(fft_d1[28]), .B(n1622), .S0(n10100), .Y(N691) );
  MX2XL U3052 ( .A(fft_d4[28]), .B(n1624), .S0(n10050), .Y(N1075) );
  MX2XL U3053 ( .A(fft_d5[28]), .B(n1718), .S0(n10030), .Y(N755) );
  MX2XL U3054 ( .A(fft_d8[28]), .B(n1720), .S0(n9980), .Y(N1139) );
  MX2XL U3055 ( .A(fft_d9[28]), .B(n1670), .S0(n9960), .Y(N723) );
  MX2XL U3056 ( .A(fft_d12[28]), .B(n1672), .S0(n9910), .Y(N1107) );
  MX2XL U3057 ( .A(fft_d13[28]), .B(n1763), .S0(n9880), .Y(N787) );
  MX2XL U3058 ( .A(fft_d1[29]), .B(n1625), .S0(n10100), .Y(N692) );
  MX2XL U3059 ( .A(fft_d4[29]), .B(n1627), .S0(n10050), .Y(N1076) );
  MX2XL U3060 ( .A(fft_d5[29]), .B(n1721), .S0(n10030), .Y(N756) );
  MX2XL U3061 ( .A(fft_d8[29]), .B(n1723), .S0(n9980), .Y(N1140) );
  MX2XL U3062 ( .A(fft_d9[29]), .B(n1673), .S0(n9960), .Y(N724) );
  MX2XL U3063 ( .A(fft_d12[29]), .B(n1675), .S0(n9910), .Y(N1108) );
  MX2XL U3064 ( .A(fft_d13[29]), .B(n1765), .S0(n9880), .Y(N788) );
  MX2XL U3065 ( .A(fft_d1[30]), .B(n1628), .S0(n10100), .Y(N693) );
  MX2XL U3066 ( .A(fft_d4[30]), .B(n1630), .S0(n10060), .Y(N1077) );
  MX2XL U3067 ( .A(fft_d5[30]), .B(n1724), .S0(n10030), .Y(N757) );
  MX2XL U3068 ( .A(fft_d8[30]), .B(n1726), .S0(n9980), .Y(N1141) );
  MX2XL U3069 ( .A(fft_d9[30]), .B(n1676), .S0(n9960), .Y(N725) );
  MX2XL U3070 ( .A(fft_d12[30]), .B(n1678), .S0(n9910), .Y(N1109) );
  MX2XL U3071 ( .A(fft_d13[30]), .B(n1767), .S0(n9880), .Y(N789) );
  MX2XL U3072 ( .A(fft_d1[31]), .B(n1631), .S0(n10100), .Y(N694) );
  MX2XL U3073 ( .A(fft_d4[31]), .B(n1633), .S0(n10060), .Y(N1078) );
  MX2XL U3074 ( .A(fft_d5[31]), .B(n1727), .S0(n10030), .Y(N758) );
  MX2XL U3075 ( .A(fft_d8[31]), .B(n1729), .S0(n9980), .Y(N1142) );
  MX2XL U3076 ( .A(fft_d9[31]), .B(n1679), .S0(n9960), .Y(N726) );
  MX2XL U3077 ( .A(fft_d12[31]), .B(n1681), .S0(n9910), .Y(N1110) );
  MX2XL U3078 ( .A(fft_d13[31]), .B(n1769), .S0(n9880), .Y(N790) );
  NOR2BX1 U3079 ( .AN(n10090), .B(n1791), .Y(N39) );
  CLKINVX3 U3080 ( .A(rst), .Y(n3149) );
  OAI221X2 U3081 ( .A0(n9800), .A1(n2855), .B0(n49), .B1(n2851), .C0(n2697), 
        .Y(stg2_real_Wn[0]) );
  NAND4X2 U3082 ( .A(n2720), .B(n2719), .C(n2718), .D(n2717), .Y(mul_2_in[14])
         );
  NAND4X2 U3083 ( .A(n2850), .B(n2849), .C(n2848), .D(n2847), .Y(mul_2_in[1])
         );
  NAND2X2 U3084 ( .A(n7300), .B(n2865), .Y(mul_0_Wn_6) );
  NAND2X2 U3085 ( .A(n197), .B(n2865), .Y(mul_0_Wn_0) );
  NAND4X2 U3086 ( .A(n2885), .B(n2884), .C(n2883), .D(n2882), .Y(mul_1_in[14])
         );
  NAND4X2 U3087 ( .A(n2897), .B(n2896), .C(n2895), .D(n2894), .Y(mul_1_in[13])
         );
  NAND4X2 U3088 ( .A(n2923), .B(n2922), .C(n2921), .D(n2920), .Y(mul_1_in[11])
         );
  NAND4X2 U3089 ( .A(n178), .B(n2948), .C(n2947), .D(n2946), .Y(mul_1_in[9])
         );
  NAND4X2 U3090 ( .A(n3053), .B(n3052), .C(n3051), .D(n3050), .Y(mul_1_in[1])
         );
  NAND4X2 U3091 ( .A(n3067), .B(n3066), .C(n3065), .D(n3064), .Y(mul_1_in[0])
         );
endmodule


module Analysis_shift_1mux_DW_cmp_0 ( A, B, GE_LT_GT_LE );
  input [31:0] A;
  input [31:0] B;
  output GE_LT_GT_LE;
  wire   n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331;

  AND2X4 U161 ( .A(n230), .B(n231), .Y(n292) );
  OAI32X4 U162 ( .A0(n251), .A1(B[30]), .A2(n295), .B0(B[31]), .B1(n250), .Y(
        n291) );
  CLKAND2X12 U163 ( .A(B[31]), .B(n250), .Y(n295) );
  NAND2BX4 U164 ( .AN(n288), .B(n298), .Y(n301) );
  OAI21X1 U165 ( .A0(n288), .A1(n289), .B0(n290), .Y(n272) );
  OAI22X1 U166 ( .A0(n291), .A1(n232), .B0(n292), .B1(n291), .Y(n290) );
  OAI22X1 U167 ( .A0(n272), .A1(n273), .B0(n274), .B1(n272), .Y(n271) );
  AOI211X2 U168 ( .A0(n255), .A1(B[24]), .B0(n299), .C0(n301), .Y(n274) );
  OAI211X2 U169 ( .A0(A[28]), .A1(n234), .B0(n294), .C0(n292), .Y(n288) );
  NAND2XL U170 ( .A(n251), .B(B[30]), .Y(n230) );
  CLKINVX1 U171 ( .A(n295), .Y(n231) );
  NAND3X1 U172 ( .A(n274), .B(n287), .C(n283), .Y(n270) );
  INVXL U173 ( .A(B[29]), .Y(n233) );
  INVX1 U174 ( .A(n287), .Y(n235) );
  AND2X2 U175 ( .A(B[27]), .B(n252), .Y(n300) );
  AND2X2 U176 ( .A(B[25]), .B(n254), .Y(n299) );
  AND2X2 U177 ( .A(B[23]), .B(n256), .Y(n281) );
  AND2X2 U178 ( .A(B[21]), .B(n258), .Y(n280) );
  AND2X2 U179 ( .A(B[19]), .B(n260), .Y(n286) );
  AND2X2 U180 ( .A(B[15]), .B(n262), .Y(n317) );
  OAI21X2 U181 ( .A0(n269), .A1(n270), .B0(n271), .Y(GE_LT_GT_LE) );
  INVXL U182 ( .A(B[17]), .Y(n238) );
  INVX1 U183 ( .A(n284), .Y(n237) );
  OAI211XL U184 ( .A0(A[16]), .A1(n239), .B0(n285), .C0(n302), .Y(n269) );
  CLKINVX1 U185 ( .A(B[12]), .Y(n242) );
  CLKINVX1 U186 ( .A(B[16]), .Y(n239) );
  CLKINVX1 U187 ( .A(B[8]), .Y(n246) );
  CLKINVX1 U188 ( .A(B[10]), .Y(n244) );
  CLKINVX1 U189 ( .A(B[9]), .Y(n245) );
  CLKINVX1 U190 ( .A(B[28]), .Y(n234) );
  CLKINVX1 U191 ( .A(B[2]), .Y(n248) );
  CLKINVX1 U192 ( .A(n279), .Y(n236) );
  CLKINVX1 U193 ( .A(n293), .Y(n232) );
  CLKINVX1 U194 ( .A(B[11]), .Y(n243) );
  CLKINVX1 U195 ( .A(n315), .Y(n240) );
  CLKINVX1 U196 ( .A(B[13]), .Y(n241) );
  CLKINVX1 U197 ( .A(B[3]), .Y(n247) );
  CLKINVX1 U198 ( .A(A[5]), .Y(n266) );
  CLKINVX1 U199 ( .A(A[0]), .Y(n249) );
  CLKINVX1 U200 ( .A(A[1]), .Y(n268) );
  CLKINVX1 U201 ( .A(A[14]), .Y(n263) );
  CLKINVX1 U202 ( .A(A[22]), .Y(n257) );
  CLKINVX1 U203 ( .A(A[15]), .Y(n262) );
  CLKINVX1 U204 ( .A(A[27]), .Y(n252) );
  CLKINVX1 U205 ( .A(A[25]), .Y(n254) );
  CLKINVX1 U206 ( .A(A[19]), .Y(n260) );
  CLKINVX1 U207 ( .A(A[7]), .Y(n264) );
  CLKINVX1 U208 ( .A(A[23]), .Y(n256) );
  CLKINVX1 U209 ( .A(A[21]), .Y(n258) );
  CLKINVX1 U210 ( .A(A[30]), .Y(n251) );
  CLKINVX1 U211 ( .A(A[31]), .Y(n250) );
  CLKINVX1 U212 ( .A(A[24]), .Y(n255) );
  CLKINVX1 U213 ( .A(A[20]), .Y(n259) );
  CLKINVX1 U214 ( .A(A[26]), .Y(n253) );
  CLKINVX1 U215 ( .A(A[18]), .Y(n261) );
  CLKINVX1 U216 ( .A(A[6]), .Y(n265) );
  CLKINVX1 U217 ( .A(A[4]), .Y(n267) );
  OAI21XL U218 ( .A0(n235), .A1(n275), .B0(n276), .Y(n273) );
  OAI22XL U219 ( .A0(n277), .A1(n278), .B0(n236), .B1(n277), .Y(n276) );
  OAI32X1 U220 ( .A0(n259), .A1(B[20]), .A2(n280), .B0(B[21]), .B1(n258), .Y(
        n278) );
  OAI32X1 U221 ( .A0(n257), .A1(B[22]), .A2(n281), .B0(B[23]), .B1(n256), .Y(
        n277) );
  OAI22XL U222 ( .A0(n282), .A1(n237), .B0(n283), .B1(n282), .Y(n275) );
  AOI32X1 U223 ( .A0(A[16]), .A1(n239), .A2(n285), .B0(n238), .B1(A[17]), .Y(
        n284) );
  OAI32X1 U224 ( .A0(n261), .A1(B[18]), .A2(n286), .B0(B[19]), .B1(n260), .Y(
        n282) );
  AOI32X1 U225 ( .A0(A[28]), .A1(n234), .A2(n294), .B0(n233), .B1(A[29]), .Y(
        n293) );
  OAI22XL U226 ( .A0(n296), .A1(n297), .B0(n298), .B1(n296), .Y(n289) );
  OAI32X1 U227 ( .A0(n255), .A1(B[24]), .A2(n299), .B0(B[25]), .B1(n254), .Y(
        n297) );
  OAI32X1 U228 ( .A0(n253), .A1(B[26]), .A2(n300), .B0(B[27]), .B1(n252), .Y(
        n296) );
  AOI21X1 U229 ( .A0(n261), .A1(B[18]), .B0(n286), .Y(n283) );
  AOI211X1 U230 ( .A0(n259), .A1(B[20]), .B0(n280), .C0(n279), .Y(n287) );
  AO21X1 U231 ( .A0(n257), .A1(B[22]), .B0(n281), .Y(n279) );
  AOI21X1 U232 ( .A0(n253), .A1(B[26]), .B0(n300), .Y(n298) );
  NAND2BX1 U233 ( .AN(A[29]), .B(B[29]), .Y(n294) );
  AOI32X1 U234 ( .A0(n303), .A1(n304), .A2(n305), .B0(n305), .B1(n306), .Y(
        n302) );
  OAI211X1 U235 ( .A0(A[8]), .A1(n246), .B0(n307), .C0(n308), .Y(n306) );
  NOR2X1 U236 ( .A(n309), .B(n310), .Y(n308) );
  OA21XL U237 ( .A0(n309), .A1(n311), .B0(n312), .Y(n305) );
  OAI22XL U238 ( .A0(n313), .A1(n240), .B0(n314), .B1(n313), .Y(n312) );
  AOI32X1 U239 ( .A0(A[12]), .A1(n242), .A2(n316), .B0(n241), .B1(A[13]), .Y(
        n315) );
  OAI32X1 U240 ( .A0(n263), .A1(B[14]), .A2(n317), .B0(B[15]), .B1(n262), .Y(
        n313) );
  AO22X1 U241 ( .A0(n318), .A1(n319), .B0(n310), .B1(n318), .Y(n311) );
  OAI21XL U242 ( .A0(A[10]), .A1(n244), .B0(n320), .Y(n310) );
  AOI32X1 U243 ( .A0(A[8]), .A1(n246), .A2(n307), .B0(n245), .B1(A[9]), .Y(
        n319) );
  NAND2BX1 U244 ( .AN(A[9]), .B(B[9]), .Y(n307) );
  AOI32X1 U245 ( .A0(A[10]), .A1(n244), .A2(n320), .B0(n243), .B1(A[11]), .Y(
        n318) );
  NAND2BX1 U246 ( .AN(A[11]), .B(B[11]), .Y(n320) );
  OAI211X1 U247 ( .A0(A[12]), .A1(n242), .B0(n316), .C0(n314), .Y(n309) );
  AOI21X1 U248 ( .A0(n263), .A1(B[14]), .B0(n317), .Y(n314) );
  NAND2BX1 U249 ( .AN(A[13]), .B(B[13]), .Y(n316) );
  OAI22XL U250 ( .A0(n321), .A1(n322), .B0(n323), .B1(n321), .Y(n304) );
  OAI32X1 U251 ( .A0(n267), .A1(B[4]), .A2(n324), .B0(B[5]), .B1(n266), .Y(
        n322) );
  OAI32X1 U252 ( .A0(n265), .A1(B[6]), .A2(n325), .B0(B[7]), .B1(n264), .Y(
        n321) );
  NAND3X1 U253 ( .A(n323), .B(n326), .C(n327), .Y(n303) );
  AOI221XL U254 ( .A0(n328), .A1(n329), .B0(B[4]), .B1(n267), .C0(n324), .Y(
        n327) );
  NOR2BX1 U255 ( .AN(B[5]), .B(A[5]), .Y(n324) );
  OAI21XL U256 ( .A0(A[2]), .A1(n248), .B0(n330), .Y(n329) );
  OAI211X1 U257 ( .A0(B[1]), .A1(n268), .B0(n331), .C0(n328), .Y(n326) );
  AOI32X1 U258 ( .A0(A[2]), .A1(n248), .A2(n330), .B0(n247), .B1(A[3]), .Y(
        n328) );
  NAND2BX1 U259 ( .AN(A[3]), .B(B[3]), .Y(n330) );
  AO22X1 U260 ( .A0(n249), .A1(B[0]), .B0(n268), .B1(B[1]), .Y(n331) );
  AOI21X1 U261 ( .A0(n265), .A1(B[6]), .B0(n325), .Y(n323) );
  AND2X1 U262 ( .A(B[7]), .B(n264), .Y(n325) );
  NAND2BX1 U263 ( .AN(A[17]), .B(B[17]), .Y(n285) );
endmodule


module Analysis_shift_1mux_DW_mult_uns_1 ( a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, b_15_, b_14_, 
        b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, 
        b_2_, b_1_, b_0_, product_31_, product_30_, product_29_, product_28_, 
        product_27_, product_26_, product_25_, product_24_, product_23_, 
        product_22_, product_21_, product_20_, product_19_, product_18_, 
        product_17_, product_16_, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_, product_2_, 
        product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_7_, a_6_, a_5_, a_4_,
         a_3_, a_2_, a_1_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_,
         b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409;

  ADDFXL U10 ( .A(n52), .B(n57), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U12 ( .A(n64), .B(n71), .CI(n12), .CO(n11), .S(product_20_) );
  ADDHXL U29 ( .A(n297), .B(n29), .CO(n28), .S(product_3_) );
  ADDFXL U31 ( .A(n194), .B(a_14_), .CI(n181), .CO(n30), .S(n31) );
  ADDFXL U32 ( .A(n182), .B(n195), .CI(n34), .CO(n32), .S(n33) );
  CMPR42X1 U33 ( .A(a_13_), .B(n208), .C(n196), .D(n183), .ICI(n37), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U34 ( .A(n209), .B(n197), .C(n184), .D(n43), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U35 ( .A(n210), .B(n185), .C(n44), .D(n48), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U36 ( .A(n221), .B(a_12_), .CI(n198), .CO(n43), .S(n44) );
  CMPR42X1 U37 ( .A(n211), .B(n53), .C(n54), .D(n49), .ICI(n50), .S(n47), 
        .ICO(n45), .CO(n46) );
  ADDFXL U38 ( .A(n199), .B(n222), .CI(n186), .CO(n48), .S(n49) );
  CMPR42X1 U39 ( .A(n200), .B(n59), .C(n55), .D(n60), .ICI(n56), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U40 ( .A(a_11_), .B(n233), .C(n223), .D(n212), .ICI(n187), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U41 ( .A(n201), .B(n68), .C(n66), .D(n61), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U42 ( .A(n213), .B(n234), .C(n224), .D(n188), .ICI(n65), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U43 ( .A(n69), .B(n76), .C(n67), .D(n74), .ICI(n70), .S(n64), .ICO(
        n62), .CO(n63) );
  CMPR42X1 U44 ( .A(n202), .B(n225), .C(n214), .D(n189), .ICI(n73), .S(n67), 
        .ICO(n65), .CO(n66) );
  ADDFXL U45 ( .A(n244), .B(a_10_), .CI(n235), .CO(n68), .S(n69) );
  CMPR42X1 U46 ( .A(n85), .B(n77), .C(n82), .D(n75), .ICI(n78), .S(n72), .ICO(
        n70), .CO(n71) );
  CMPR42X1 U47 ( .A(n236), .B(n215), .C(n226), .D(n84), .ICI(n81), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U48 ( .A(n203), .B(n245), .CI(n190), .CO(n76), .S(n77) );
  CMPR42X1 U49 ( .A(n86), .B(n94), .C(n91), .D(n83), .ICI(n87), .S(n80), .ICO(
        n78), .CO(n79) );
  CMPR42X1 U50 ( .A(n237), .B(n216), .C(n227), .D(n90), .ICI(n93), .S(n83), 
        .ICO(n81), .CO(n82) );
  CMPR42X1 U51 ( .A(a_9_), .B(n254), .C(n246), .D(n204), .ICI(n191), .S(n86), 
        .ICO(n84), .CO(n85) );
  CMPR42X1 U52 ( .A(n103), .B(n95), .C(n92), .D(n100), .ICI(n96), .S(n89), 
        .ICO(n87), .CO(n88) );
  CMPR42X1 U53 ( .A(n255), .B(n238), .C(n247), .D(n99), .ICI(n102), .S(n92), 
        .ICO(n90), .CO(n91) );
  CMPR42X1 U54 ( .A(n217), .B(n205), .C(n228), .D(n192), .ICI(b_8_), .S(n95), 
        .ICO(n93), .CO(n94) );
  CMPR42X1 U55 ( .A(n113), .B(n104), .C(n111), .D(n107), .ICI(n101), .S(n98), 
        .ICO(n96), .CO(n97) );
  CMPR42X1 U56 ( .A(n239), .B(n218), .C(n229), .D(n106), .ICI(n110), .S(n101), 
        .ICO(n99), .CO(n100) );
  CMPR42X1 U57 ( .A(n256), .B(n206), .C(n248), .D(n193), .ICI(n115), .S(n104), 
        .ICO(n102), .CO(n103) );
  CMPR42X1 U60 ( .A(n123), .B(n114), .C(n121), .D(n112), .ICI(n117), .S(n109), 
        .ICO(n107), .CO(n108) );
  CMPR42X1 U61 ( .A(n249), .B(n230), .C(n125), .D(n120), .ICI(n116), .S(n112), 
        .ICO(n110), .CO(n111) );
  ADDFXL U62 ( .A(n264), .B(n240), .CI(n257), .CO(n113), .S(n114) );
  ADDHXL U63 ( .A(n219), .B(n207), .CO(n115), .S(n116) );
  CMPR42X1 U64 ( .A(n126), .B(n131), .C(n124), .D(n122), .ICI(n127), .S(n119), 
        .ICO(n117), .CO(n118) );
  CMPR42X1 U65 ( .A(n250), .B(n265), .C(n258), .D(n133), .ICI(n130), .S(n122), 
        .ICO(n120), .CO(n121) );
  ADDFXL U66 ( .A(n220), .B(n271), .CI(n241), .CO(n123), .S(n124) );
  ADDHXL U67 ( .A(a_7_), .B(n231), .CO(n125), .S(n126) );
  CMPR42X1 U68 ( .A(n141), .B(n134), .C(n139), .D(n132), .ICI(n135), .S(n129), 
        .ICO(n127), .CO(n128) );
  CMPR42X1 U69 ( .A(n272), .B(n251), .C(n266), .D(n259), .ICI(n138), .S(n132), 
        .ICO(n130), .CO(n131) );
  ADDHXL U70 ( .A(n242), .B(n232), .CO(n133), .S(n134) );
  CMPR42X1 U71 ( .A(n267), .B(n142), .C(n146), .D(n140), .ICI(n143), .S(n137), 
        .ICO(n135), .CO(n136) );
  CMPR42X1 U72 ( .A(n278), .B(n243), .C(n273), .D(n260), .ICI(n148), .S(n140), 
        .ICO(n138), .CO(n139) );
  ADDHXL U73 ( .A(a_6_), .B(n252), .CO(n141), .S(n142) );
  CMPR42X1 U74 ( .A(n155), .B(n149), .C(n153), .D(n150), .ICI(n147), .S(n145), 
        .ICO(n143), .CO(n144) );
  ADDFXL U75 ( .A(n274), .B(n268), .CI(n279), .CO(n146), .S(n147) );
  ADDHXL U76 ( .A(n261), .B(n253), .CO(n148), .S(n149) );
  ADDFXL U78 ( .A(n262), .B(n284), .CI(n275), .CO(n153), .S(n154) );
  CMPR42X1 U80 ( .A(n285), .B(n281), .C(n165), .D(n162), .ICI(n161), .S(n159), 
        .ICO(n157), .CO(n158) );
  ADDHXL U81 ( .A(n276), .B(n270), .CO(n160), .S(n161) );
  CMPR42X1 U82 ( .A(n289), .B(n277), .C(n286), .D(n169), .ICI(n166), .S(n164), 
        .ICO(n162), .CO(n163) );
  ADDFXL U84 ( .A(n173), .B(n287), .CI(n170), .CO(n167), .S(n168) );
  ADDHXL U85 ( .A(n290), .B(n283), .CO(n169), .S(n170) );
  ADDFXL U86 ( .A(n288), .B(n291), .CI(n175), .CO(n171), .S(n172) );
  ADDHXL U87 ( .A(a_3_), .B(n293), .CO(n173), .S(n174) );
  ADDFHX2 U243 ( .A(n88), .B(n80), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFHX4 U244 ( .A(n179), .B(a_15_), .CI(n2), .CO(n1), .S(product_30_) );
  BUFX16 U245 ( .A(n406), .Y(n392) );
  CLKINVX12 U246 ( .A(b_3_), .Y(n406) );
  CMPR42X2 U247 ( .A(n280), .B(n160), .C(n156), .D(n157), .ICI(n154), .S(n152), 
        .ICO(n150), .CO(n151) );
  ADDHX1 U248 ( .A(a_5_), .B(n269), .CO(n155), .S(n156) );
  NOR2XL U249 ( .A(n391), .B(n381), .Y(n203) );
  NOR2XL U250 ( .A(n391), .B(n382), .Y(n216) );
  NOR2XL U251 ( .A(n391), .B(n384), .Y(n239) );
  NOR2XL U252 ( .A(n391), .B(n385), .Y(n249) );
  NOR2XL U253 ( .A(n391), .B(n386), .Y(n258) );
  NOR2XL U254 ( .A(n387), .B(n391), .Y(n266) );
  NOR2XL U255 ( .A(n391), .B(n388), .Y(n273) );
  NOR2XL U256 ( .A(n392), .B(n391), .Y(n289) );
  NOR2XL U257 ( .A(n407), .B(n391), .Y(n290) );
  NOR2XL U258 ( .A(n394), .B(n391), .Y(n292) );
  NOR2X4 U259 ( .A(n393), .B(n391), .Y(n291) );
  NOR2X2 U260 ( .A(n394), .B(n390), .Y(n288) );
  NOR2X2 U261 ( .A(n393), .B(n390), .Y(n287) );
  NOR2XL U262 ( .A(n391), .B(n390), .Y(n284) );
  NOR2XL U263 ( .A(n407), .B(n390), .Y(n286) );
  NOR2XL U264 ( .A(n392), .B(n390), .Y(n285) );
  BUFX8 U265 ( .A(n404), .Y(n390) );
  NOR2X2 U266 ( .A(n394), .B(n389), .Y(n283) );
  NOR2XL U267 ( .A(n393), .B(n389), .Y(n282) );
  NOR2XL U268 ( .A(n407), .B(n389), .Y(n281) );
  NOR2XL U269 ( .A(n390), .B(n389), .Y(n278) );
  NOR2XL U270 ( .A(n392), .B(n389), .Y(n280) );
  NOR2XL U271 ( .A(n391), .B(n389), .Y(n279) );
  BUFX12 U272 ( .A(n403), .Y(n389) );
  ADDFHX4 U273 ( .A(n159), .B(n163), .CI(n23), .CO(n22), .S(product_9_) );
  NOR2X8 U274 ( .A(n394), .B(n393), .Y(n298) );
  NOR2X4 U275 ( .A(n393), .B(n407), .Y(n296) );
  NOR2X2 U276 ( .A(n393), .B(n392), .Y(n294) );
  BUFX12 U277 ( .A(n408), .Y(n393) );
  NOR2X2 U278 ( .A(n407), .B(n392), .Y(n293) );
  INVX20 U279 ( .A(b_5_), .Y(n404) );
  ADDHX1 U280 ( .A(n294), .B(n292), .CO(n175), .S(n176) );
  INVX20 U281 ( .A(b_2_), .Y(n407) );
  ADDHX2 U282 ( .A(a_2_), .B(n296), .CO(n177), .S(n178) );
  CLKBUFX3 U283 ( .A(n401), .Y(n387) );
  CLKBUFX3 U284 ( .A(n402), .Y(n388) );
  CLKBUFX3 U285 ( .A(n400), .Y(n386) );
  CLKBUFX3 U286 ( .A(n399), .Y(n385) );
  CLKBUFX3 U287 ( .A(n397), .Y(n383) );
  CLKBUFX3 U288 ( .A(n396), .Y(n382) );
  CLKBUFX3 U289 ( .A(n398), .Y(n384) );
  CLKBUFX3 U290 ( .A(n395), .Y(n381) );
  CLKINVX1 U291 ( .A(b_1_), .Y(n408) );
  CLKBUFX8 U292 ( .A(n409), .Y(n394) );
  ADDFX2 U293 ( .A(n72), .B(n79), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFX2 U294 ( .A(n58), .B(n63), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U295 ( .A(n47), .B(n51), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U296 ( .A(n39), .B(n41), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U297 ( .A(n33), .B(n35), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U298 ( .A(n42), .B(n46), .CI(n8), .CO(n7), .S(product_24_) );
  CLKINVX1 U299 ( .A(n1), .Y(product_31_) );
  CLKINVX1 U300 ( .A(b_0_), .Y(n409) );
  ADDHX1 U301 ( .A(a_1_), .B(n298), .CO(n29), .S(product_2_) );
  NAND2XL U302 ( .A(b_15_), .B(b_14_), .Y(n179) );
  NAND2XL U303 ( .A(b_15_), .B(b_13_), .Y(n180) );
  NAND2XL U304 ( .A(b_8_), .B(n388), .Y(n106) );
  NAND2XL U305 ( .A(b_15_), .B(b_3_), .Y(n190) );
  ADDFHX4 U306 ( .A(n145), .B(n151), .CI(n21), .CO(n20), .S(product_11_) );
  ADDHX1 U307 ( .A(a_4_), .B(n282), .CO(n165), .S(n166) );
  ADDFHX2 U308 ( .A(n167), .B(n164), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFHX2 U309 ( .A(n109), .B(n118), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFHX2 U310 ( .A(n89), .B(n97), .CI(n15), .CO(n14), .S(product_17_) );
  ADDFX1 U311 ( .A(n119), .B(n128), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFX1 U312 ( .A(n137), .B(n144), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFX1 U313 ( .A(n129), .B(n136), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFX1 U314 ( .A(n98), .B(n108), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFX2 U315 ( .A(n172), .B(n174), .CI(n26), .CO(n25), .S(product_6_) );
  BUFX4 U316 ( .A(n405), .Y(n391) );
  ADDFX1 U317 ( .A(n168), .B(n171), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFX1 U318 ( .A(n152), .B(n158), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFX1 U319 ( .A(n178), .B(n295), .CI(n28), .CO(n27), .S(product_4_) );
  ADDFX1 U320 ( .A(n176), .B(n177), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFHX1 U321 ( .A(n30), .B(n180), .CI(n3), .CO(n2), .S(product_29_) );
  NOR2XL U322 ( .A(n387), .B(n393), .Y(n269) );
  NOR2XL U323 ( .A(n393), .B(n385), .Y(n252) );
  NOR2XL U324 ( .A(n393), .B(n383), .Y(n231) );
  NOR2XL U325 ( .A(n391), .B(n383), .Y(n228) );
  NAND2XL U326 ( .A(b_15_), .B(b_1_), .Y(n192) );
  NOR2XL U327 ( .A(n407), .B(n381), .Y(n205) );
  NOR2XL U328 ( .A(n390), .B(n385), .Y(n248) );
  NAND2XL U329 ( .A(b_15_), .B(b_0_), .Y(n193) );
  NOR2XL U330 ( .A(n393), .B(n381), .Y(n206) );
  NOR2XL U331 ( .A(n387), .B(n384), .Y(n235) );
  NOR2XL U332 ( .A(n386), .B(n385), .Y(n244) );
  NOR2XL U333 ( .A(n387), .B(n381), .Y(n199) );
  NAND2XL U334 ( .A(b_15_), .B(b_7_), .Y(n186) );
  NOR2XL U335 ( .A(n385), .B(n383), .Y(n222) );
  NAND2XL U336 ( .A(b_15_), .B(b_2_), .Y(n191) );
  NOR2XL U337 ( .A(n392), .B(n381), .Y(n204) );
  NOR2XL U338 ( .A(n388), .B(n385), .Y(n246) );
  NAND2XL U339 ( .A(b_15_), .B(b_6_), .Y(n187) );
  NOR2XL U340 ( .A(n387), .B(n382), .Y(n212) );
  NOR2XL U341 ( .A(n386), .B(n383), .Y(n223) );
  NOR2XL U342 ( .A(n389), .B(n382), .Y(n214) );
  NAND2XL U343 ( .A(b_15_), .B(b_4_), .Y(n189) );
  NOR2XL U344 ( .A(n388), .B(n383), .Y(n225) );
  NOR2XL U345 ( .A(n387), .B(n383), .Y(n224) );
  NAND2XL U346 ( .A(b_15_), .B(b_5_), .Y(n188) );
  NOR2XL U347 ( .A(n386), .B(n384), .Y(n234) );
  NOR2XL U348 ( .A(n386), .B(n381), .Y(n198) );
  NOR2XL U349 ( .A(n384), .B(n383), .Y(n221) );
  NOR2XL U350 ( .A(n385), .B(n382), .Y(n210) );
  NAND2XL U351 ( .A(b_15_), .B(b_8_), .Y(n185) );
  NAND2XL U352 ( .A(b_15_), .B(b_9_), .Y(n184) );
  NOR2XL U353 ( .A(n385), .B(n381), .Y(n197) );
  NOR2XL U354 ( .A(n384), .B(n382), .Y(n209) );
  NOR2XL U355 ( .A(n382), .B(n381), .Y(n194) );
  NAND2XL U356 ( .A(b_15_), .B(b_12_), .Y(n181) );
  NAND2XL U357 ( .A(b_15_), .B(b_11_), .Y(n182) );
  NOR2XL U358 ( .A(n383), .B(n381), .Y(n195) );
  NOR2XL U359 ( .A(n384), .B(n381), .Y(n196) );
  NAND2XL U360 ( .A(b_15_), .B(b_10_), .Y(n183) );
  NOR2XL U361 ( .A(n383), .B(n382), .Y(n208) );
  ADDFXL U362 ( .A(n38), .B(n36), .CI(n6), .CO(n5), .S(product_26_) );
  ADDFXL U363 ( .A(n32), .B(n31), .CI(n4), .CO(n3), .S(product_28_) );
  INVXL U364 ( .A(b_4_), .Y(n405) );
  INVXL U365 ( .A(b_6_), .Y(n403) );
  INVXL U366 ( .A(b_8_), .Y(n401) );
  INVXL U367 ( .A(b_13_), .Y(n396) );
  INVXL U368 ( .A(b_11_), .Y(n398) );
  INVXL U369 ( .A(b_7_), .Y(n402) );
  INVXL U370 ( .A(b_9_), .Y(n400) );
  INVXL U371 ( .A(b_10_), .Y(n399) );
  INVXL U372 ( .A(b_12_), .Y(n397) );
  INVXL U373 ( .A(b_14_), .Y(n395) );
  CLKBUFX2 U374 ( .A(b_0_), .Y(product_0_) );
  NOR2X1 U375 ( .A(n394), .B(n407), .Y(n297) );
  NOR2X1 U376 ( .A(n394), .B(n392), .Y(n295) );
  NOR2X1 U377 ( .A(n394), .B(n388), .Y(n277) );
  NOR2X1 U378 ( .A(n393), .B(n388), .Y(n276) );
  NOR2X1 U379 ( .A(n407), .B(n388), .Y(n275) );
  NOR2X1 U380 ( .A(n392), .B(n388), .Y(n274) );
  NOR2X1 U381 ( .A(n390), .B(n388), .Y(n272) );
  NOR2X1 U382 ( .A(n389), .B(n388), .Y(n271) );
  NOR2X1 U383 ( .A(n387), .B(n394), .Y(n270) );
  NOR2X1 U384 ( .A(n387), .B(n407), .Y(n268) );
  NOR2X1 U385 ( .A(n387), .B(n392), .Y(n267) );
  NOR2X1 U386 ( .A(n387), .B(n390), .Y(n265) );
  NOR2X1 U387 ( .A(n387), .B(n389), .Y(n264) );
  NOR2X1 U388 ( .A(n394), .B(n386), .Y(n262) );
  NOR2X1 U389 ( .A(n393), .B(n386), .Y(n261) );
  NOR2X1 U390 ( .A(n407), .B(n386), .Y(n260) );
  NOR2X1 U391 ( .A(n392), .B(n386), .Y(n259) );
  NOR2X1 U392 ( .A(n390), .B(n386), .Y(n257) );
  NOR2X1 U393 ( .A(n389), .B(n386), .Y(n256) );
  NOR2X1 U394 ( .A(n388), .B(n386), .Y(n255) );
  NOR2X1 U395 ( .A(n387), .B(n386), .Y(n254) );
  NOR2X1 U396 ( .A(n394), .B(n385), .Y(n253) );
  NOR2X1 U397 ( .A(n407), .B(n385), .Y(n251) );
  NOR2X1 U398 ( .A(n392), .B(n385), .Y(n250) );
  NOR2X1 U399 ( .A(n389), .B(n385), .Y(n247) );
  NOR2X1 U400 ( .A(n387), .B(n385), .Y(n245) );
  NOR2X1 U401 ( .A(n394), .B(n384), .Y(n243) );
  NOR2X1 U402 ( .A(n393), .B(n384), .Y(n242) );
  NOR2X1 U403 ( .A(n407), .B(n384), .Y(n241) );
  NOR2X1 U404 ( .A(n392), .B(n384), .Y(n240) );
  NOR2X1 U405 ( .A(n390), .B(n384), .Y(n238) );
  NOR2X1 U406 ( .A(n389), .B(n384), .Y(n237) );
  NOR2X1 U407 ( .A(n388), .B(n384), .Y(n236) );
  NOR2X1 U408 ( .A(n385), .B(n384), .Y(n233) );
  NOR2X1 U409 ( .A(n394), .B(n383), .Y(n232) );
  NOR2X1 U410 ( .A(n407), .B(n383), .Y(n230) );
  NOR2X1 U411 ( .A(n392), .B(n383), .Y(n229) );
  NOR2X1 U412 ( .A(n390), .B(n383), .Y(n227) );
  NOR2X1 U413 ( .A(n389), .B(n383), .Y(n226) );
  NOR2X1 U414 ( .A(n394), .B(n382), .Y(n220) );
  NOR2X1 U415 ( .A(n393), .B(n382), .Y(n219) );
  NOR2X1 U416 ( .A(n407), .B(n382), .Y(n218) );
  NOR2X1 U417 ( .A(n392), .B(n382), .Y(n217) );
  NOR2X1 U418 ( .A(n390), .B(n382), .Y(n215) );
  NOR2X1 U419 ( .A(n388), .B(n382), .Y(n213) );
  NOR2X1 U420 ( .A(n386), .B(n382), .Y(n211) );
  NOR2X1 U421 ( .A(n394), .B(n381), .Y(n207) );
  NOR2X1 U422 ( .A(n390), .B(n381), .Y(n202) );
  NOR2X1 U423 ( .A(n389), .B(n381), .Y(n201) );
  NOR2X1 U424 ( .A(n388), .B(n381), .Y(n200) );
endmodule


module Analysis_shift_1mux_DW_mult_uns_0 ( a_15_, a_14_, a_13_, a_12_, a_11_, 
        a_10_, a_9_, a_7_, a_6_, a_5_, a_4_, a_3_, a_2_, a_1_, b_15_, b_14_, 
        b_13_, b_12_, b_11_, b_10_, b_9_, b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, 
        b_2_, b_1_, b_0_, product_31_, product_30_, product_29_, product_28_, 
        product_27_, product_26_, product_25_, product_24_, product_23_, 
        product_22_, product_21_, product_20_, product_19_, product_18_, 
        product_17_, product_16_, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_, product_2_, 
        product_0_ );
  input a_15_, a_14_, a_13_, a_12_, a_11_, a_10_, a_9_, a_7_, a_6_, a_5_, a_4_,
         a_3_, a_2_, a_1_, b_15_, b_14_, b_13_, b_12_, b_11_, b_10_, b_9_,
         b_8_, b_7_, b_6_, b_5_, b_4_, b_3_, b_2_, b_1_, b_0_;
  output product_31_, product_30_, product_29_, product_28_, product_27_,
         product_26_, product_25_, product_24_, product_23_, product_22_,
         product_21_, product_20_, product_19_, product_18_, product_17_,
         product_16_, product_15_, product_14_, product_13_, product_12_,
         product_11_, product_10_, product_9_, product_8_, product_7_,
         product_6_, product_5_, product_4_, product_3_, product_2_,
         product_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407;

  ADDFXL U10 ( .A(n52), .B(n57), .CI(n10), .CO(n9), .S(product_22_) );
  ADDFXL U12 ( .A(n64), .B(n71), .CI(n12), .CO(n11), .S(product_20_) );
  ADDHXL U29 ( .A(n297), .B(n29), .CO(n28), .S(product_3_) );
  ADDFXL U31 ( .A(n194), .B(a_14_), .CI(n181), .CO(n30), .S(n31) );
  ADDFXL U32 ( .A(n182), .B(n195), .CI(n34), .CO(n32), .S(n33) );
  CMPR42X1 U33 ( .A(a_13_), .B(n208), .C(n196), .D(n183), .ICI(n37), .S(n36), 
        .ICO(n34), .CO(n35) );
  CMPR42X1 U34 ( .A(n209), .B(n197), .C(n184), .D(n43), .ICI(n40), .S(n39), 
        .ICO(n37), .CO(n38) );
  CMPR42X1 U35 ( .A(n210), .B(n185), .C(n44), .D(n48), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U36 ( .A(n221), .B(a_12_), .CI(n198), .CO(n43), .S(n44) );
  CMPR42X1 U37 ( .A(n211), .B(n53), .C(n54), .D(n49), .ICI(n50), .S(n47), 
        .ICO(n45), .CO(n46) );
  ADDFXL U38 ( .A(n199), .B(n222), .CI(n186), .CO(n48), .S(n49) );
  CMPR42X1 U39 ( .A(n200), .B(n59), .C(n55), .D(n60), .ICI(n56), .S(n52), 
        .ICO(n50), .CO(n51) );
  CMPR42X1 U40 ( .A(a_11_), .B(n233), .C(n223), .D(n212), .ICI(n187), .S(n55), 
        .ICO(n53), .CO(n54) );
  CMPR42X1 U41 ( .A(n201), .B(n68), .C(n66), .D(n61), .ICI(n62), .S(n58), 
        .ICO(n56), .CO(n57) );
  CMPR42X1 U42 ( .A(n213), .B(n234), .C(n224), .D(n188), .ICI(n65), .S(n61), 
        .ICO(n59), .CO(n60) );
  CMPR42X1 U43 ( .A(n69), .B(n76), .C(n67), .D(n74), .ICI(n70), .S(n64), .ICO(
        n62), .CO(n63) );
  CMPR42X1 U44 ( .A(n202), .B(n225), .C(n214), .D(n189), .ICI(n73), .S(n67), 
        .ICO(n65), .CO(n66) );
  ADDFXL U45 ( .A(n244), .B(a_10_), .CI(n235), .CO(n68), .S(n69) );
  CMPR42X1 U46 ( .A(n85), .B(n77), .C(n82), .D(n75), .ICI(n78), .S(n72), .ICO(
        n70), .CO(n71) );
  CMPR42X1 U47 ( .A(n236), .B(n215), .C(n226), .D(n84), .ICI(n81), .S(n75), 
        .ICO(n73), .CO(n74) );
  ADDFXL U48 ( .A(n203), .B(n245), .CI(n190), .CO(n76), .S(n77) );
  CMPR42X1 U49 ( .A(n86), .B(n94), .C(n91), .D(n83), .ICI(n87), .S(n80), .ICO(
        n78), .CO(n79) );
  CMPR42X1 U50 ( .A(n237), .B(n216), .C(n227), .D(n90), .ICI(n93), .S(n83), 
        .ICO(n81), .CO(n82) );
  CMPR42X1 U51 ( .A(a_9_), .B(n254), .C(n246), .D(n204), .ICI(n191), .S(n86), 
        .ICO(n84), .CO(n85) );
  CMPR42X1 U52 ( .A(n103), .B(n95), .C(n92), .D(n100), .ICI(n96), .S(n89), 
        .ICO(n87), .CO(n88) );
  CMPR42X1 U53 ( .A(n255), .B(n238), .C(n247), .D(n99), .ICI(n102), .S(n92), 
        .ICO(n90), .CO(n91) );
  CMPR42X1 U54 ( .A(n217), .B(n205), .C(n228), .D(n192), .ICI(b_8_), .S(n95), 
        .ICO(n93), .CO(n94) );
  CMPR42X1 U55 ( .A(n113), .B(n104), .C(n111), .D(n107), .ICI(n101), .S(n98), 
        .ICO(n96), .CO(n97) );
  CMPR42X1 U56 ( .A(n239), .B(n218), .C(n229), .D(n106), .ICI(n110), .S(n101), 
        .ICO(n99), .CO(n100) );
  CMPR42X1 U57 ( .A(n256), .B(n206), .C(n248), .D(n193), .ICI(n115), .S(n104), 
        .ICO(n102), .CO(n103) );
  CMPR42X1 U60 ( .A(n123), .B(n114), .C(n121), .D(n112), .ICI(n117), .S(n109), 
        .ICO(n107), .CO(n108) );
  CMPR42X1 U61 ( .A(n249), .B(n230), .C(n125), .D(n120), .ICI(n116), .S(n112), 
        .ICO(n110), .CO(n111) );
  ADDFXL U62 ( .A(n264), .B(n240), .CI(n257), .CO(n113), .S(n114) );
  ADDHXL U63 ( .A(n219), .B(n207), .CO(n115), .S(n116) );
  CMPR42X1 U64 ( .A(n126), .B(n131), .C(n124), .D(n122), .ICI(n127), .S(n119), 
        .ICO(n117), .CO(n118) );
  CMPR42X1 U65 ( .A(n250), .B(n265), .C(n258), .D(n133), .ICI(n130), .S(n122), 
        .ICO(n120), .CO(n121) );
  ADDFXL U66 ( .A(n220), .B(n271), .CI(n241), .CO(n123), .S(n124) );
  ADDHXL U67 ( .A(a_7_), .B(n231), .CO(n125), .S(n126) );
  CMPR42X1 U68 ( .A(n141), .B(n134), .C(n139), .D(n132), .ICI(n135), .S(n129), 
        .ICO(n127), .CO(n128) );
  CMPR42X1 U69 ( .A(n272), .B(n251), .C(n266), .D(n259), .ICI(n138), .S(n132), 
        .ICO(n130), .CO(n131) );
  ADDHXL U70 ( .A(n242), .B(n232), .CO(n133), .S(n134) );
  CMPR42X1 U72 ( .A(n278), .B(n243), .C(n273), .D(n260), .ICI(n148), .S(n140), 
        .ICO(n138), .CO(n139) );
  ADDFXL U75 ( .A(n274), .B(n268), .CI(n279), .CO(n146), .S(n147) );
  CMPR42X1 U77 ( .A(n280), .B(n160), .C(n156), .D(n157), .ICI(n154), .S(n152), 
        .ICO(n150), .CO(n151) );
  ADDFXL U78 ( .A(n262), .B(n284), .CI(n275), .CO(n153), .S(n154) );
  CMPR42X1 U80 ( .A(n285), .B(n281), .C(n165), .D(n162), .ICI(n161), .S(n159), 
        .ICO(n157), .CO(n158) );
  ADDHXL U81 ( .A(n276), .B(n270), .CO(n160), .S(n161) );
  CMPR42X1 U82 ( .A(n289), .B(n277), .C(n286), .D(n169), .ICI(n166), .S(n164), 
        .ICO(n162), .CO(n163) );
  ADDFXL U84 ( .A(n173), .B(n287), .CI(n170), .CO(n167), .S(n168) );
  ADDHXL U85 ( .A(n290), .B(n283), .CO(n169), .S(n170) );
  ADDFXL U86 ( .A(n288), .B(n291), .CI(n175), .CO(n171), .S(n172) );
  ADDHXL U88 ( .A(n294), .B(n292), .CO(n175), .S(n176) );
  NOR2XL U243 ( .A(n387), .B(n392), .Y(n270) );
  NOR2XL U244 ( .A(n387), .B(n405), .Y(n268) );
  BUFX4 U245 ( .A(n399), .Y(n387) );
  CMPR42X2 U246 ( .A(n267), .B(n142), .C(n146), .D(n140), .ICI(n143), .S(n137), 
        .ICO(n135), .CO(n136) );
  ADDHX1 U247 ( .A(a_6_), .B(n252), .CO(n141), .S(n142) );
  CMPR42X2 U248 ( .A(n155), .B(n149), .C(n153), .D(n150), .ICI(n147), .S(n145), 
        .ICO(n143), .CO(n144) );
  ADDHX2 U249 ( .A(n261), .B(n253), .CO(n148), .S(n149) );
  ADDFHX4 U250 ( .A(n152), .B(n158), .CI(n22), .CO(n21), .S(product_10_) );
  ADDFHX1 U251 ( .A(n159), .B(n163), .CI(n23), .CO(n22), .S(product_9_) );
  CLKINVX16 U252 ( .A(b_0_), .Y(n407) );
  ADDFHX2 U253 ( .A(n179), .B(a_15_), .CI(n2), .CO(n1), .S(product_30_) );
  BUFX20 U254 ( .A(n403), .Y(n390) );
  INVX20 U255 ( .A(b_4_), .Y(n403) );
  BUFX20 U256 ( .A(n402), .Y(n389) );
  INVX20 U257 ( .A(b_5_), .Y(n402) );
  NOR2X2 U258 ( .A(n392), .B(n390), .Y(n292) );
  NOR2X2 U259 ( .A(n406), .B(n390), .Y(n291) );
  NOR2X2 U260 ( .A(n405), .B(n390), .Y(n290) );
  NOR2X2 U261 ( .A(n391), .B(n390), .Y(n289) );
  NOR2XL U262 ( .A(n390), .B(n389), .Y(n284) );
  NOR2XL U263 ( .A(n390), .B(n388), .Y(n273) );
  NOR2XL U264 ( .A(n389), .B(n388), .Y(n272) );
  BUFX12 U265 ( .A(n400), .Y(n388) );
  NOR2X2 U266 ( .A(n392), .B(n406), .Y(n298) );
  NOR2X4 U267 ( .A(n406), .B(n405), .Y(n296) );
  NOR2X4 U268 ( .A(n406), .B(n391), .Y(n294) );
  NOR2X1 U269 ( .A(n406), .B(n401), .Y(n282) );
  INVX8 U270 ( .A(b_1_), .Y(n406) );
  NOR2XL U271 ( .A(n392), .B(n391), .Y(n295) );
  NOR2X2 U272 ( .A(n405), .B(n391), .Y(n293) );
  NOR2X2 U273 ( .A(n391), .B(n389), .Y(n285) );
  BUFX20 U274 ( .A(n404), .Y(n391) );
  INVX20 U275 ( .A(b_6_), .Y(n401) );
  NOR2XL U276 ( .A(n391), .B(n383), .Y(n229) );
  NOR2XL U277 ( .A(n391), .B(n382), .Y(n217) );
  NOR2XL U278 ( .A(n391), .B(n384), .Y(n240) );
  NOR2XL U279 ( .A(n391), .B(n385), .Y(n250) );
  NOR2XL U280 ( .A(n387), .B(n391), .Y(n267) );
  NOR2XL U281 ( .A(n391), .B(n386), .Y(n259) );
  NOR2XL U282 ( .A(n391), .B(n401), .Y(n280) );
  NOR2XL U283 ( .A(n391), .B(n388), .Y(n274) );
  NOR2X2 U284 ( .A(n405), .B(n389), .Y(n286) );
  CLKINVX20 U285 ( .A(b_2_), .Y(n405) );
  CMPR22X2 U286 ( .A(a_2_), .B(n296), .CO(n177), .S(n178) );
  INVX16 U287 ( .A(b_3_), .Y(n404) );
  ADDHX2 U288 ( .A(a_3_), .B(n293), .CO(n173), .S(n174) );
  CLKBUFX3 U289 ( .A(n398), .Y(n386) );
  CLKBUFX3 U290 ( .A(n397), .Y(n385) );
  CLKBUFX3 U291 ( .A(n395), .Y(n383) );
  CLKBUFX3 U292 ( .A(n394), .Y(n382) );
  CLKBUFX3 U293 ( .A(n396), .Y(n384) );
  CLKBUFX3 U294 ( .A(n393), .Y(n381) );
  BUFX6 U295 ( .A(n407), .Y(n392) );
  ADDFXL U296 ( .A(n72), .B(n79), .CI(n13), .CO(n12), .S(product_19_) );
  ADDFXL U297 ( .A(n58), .B(n63), .CI(n11), .CO(n10), .S(product_21_) );
  ADDFXL U298 ( .A(n47), .B(n51), .CI(n9), .CO(n8), .S(product_23_) );
  ADDFXL U299 ( .A(n39), .B(n41), .CI(n7), .CO(n6), .S(product_25_) );
  ADDFXL U300 ( .A(n33), .B(n35), .CI(n5), .CO(n4), .S(product_27_) );
  ADDFXL U301 ( .A(n88), .B(n80), .CI(n14), .CO(n13), .S(product_18_) );
  ADDFXL U302 ( .A(n42), .B(n46), .CI(n8), .CO(n7), .S(product_24_) );
  ADDHX2 U303 ( .A(a_1_), .B(n298), .CO(n29), .S(product_2_) );
  NAND2XL U304 ( .A(b_15_), .B(b_14_), .Y(n179) );
  NAND2XL U305 ( .A(b_15_), .B(b_13_), .Y(n180) );
  NAND2XL U306 ( .A(b_8_), .B(n388), .Y(n106) );
  NAND2XL U307 ( .A(b_15_), .B(b_3_), .Y(n190) );
  ADDFHX2 U308 ( .A(n89), .B(n97), .CI(n15), .CO(n14), .S(product_17_) );
  ADDHX1 U309 ( .A(a_5_), .B(n269), .CO(n155), .S(n156) );
  ADDFHX4 U310 ( .A(n145), .B(n151), .CI(n21), .CO(n20), .S(product_11_) );
  ADDHX1 U311 ( .A(a_4_), .B(n282), .CO(n165), .S(n166) );
  ADDFHX2 U312 ( .A(n167), .B(n164), .CI(n24), .CO(n23), .S(product_8_) );
  ADDFHX2 U313 ( .A(n109), .B(n118), .CI(n17), .CO(n16), .S(product_15_) );
  ADDFX1 U314 ( .A(n119), .B(n128), .CI(n18), .CO(n17), .S(product_14_) );
  ADDFX1 U315 ( .A(n137), .B(n144), .CI(n20), .CO(n19), .S(product_12_) );
  ADDFX1 U316 ( .A(n129), .B(n136), .CI(n19), .CO(n18), .S(product_13_) );
  ADDFX1 U317 ( .A(n98), .B(n108), .CI(n16), .CO(n15), .S(product_16_) );
  ADDFX2 U318 ( .A(n172), .B(n174), .CI(n26), .CO(n25), .S(product_6_) );
  ADDFX1 U319 ( .A(n168), .B(n171), .CI(n25), .CO(n24), .S(product_7_) );
  ADDFX1 U320 ( .A(n178), .B(n295), .CI(n28), .CO(n27), .S(product_4_) );
  ADDFX1 U321 ( .A(n176), .B(n177), .CI(n27), .CO(n26), .S(product_5_) );
  ADDFHX1 U322 ( .A(n30), .B(n180), .CI(n3), .CO(n2), .S(product_29_) );
  NOR2XL U323 ( .A(n387), .B(n406), .Y(n269) );
  NOR2XL U324 ( .A(n406), .B(n385), .Y(n252) );
  NOR2XL U325 ( .A(n406), .B(n383), .Y(n231) );
  NOR2XL U326 ( .A(n390), .B(n383), .Y(n228) );
  NAND2XL U327 ( .A(b_15_), .B(b_1_), .Y(n192) );
  NOR2XL U328 ( .A(n405), .B(n381), .Y(n205) );
  NOR2XL U329 ( .A(n389), .B(n385), .Y(n248) );
  NAND2XL U330 ( .A(b_15_), .B(b_0_), .Y(n193) );
  NOR2XL U331 ( .A(n406), .B(n381), .Y(n206) );
  NOR2XL U332 ( .A(n387), .B(n384), .Y(n235) );
  NOR2XL U333 ( .A(n386), .B(n385), .Y(n244) );
  NOR2XL U334 ( .A(n387), .B(n381), .Y(n199) );
  NAND2XL U335 ( .A(b_15_), .B(b_7_), .Y(n186) );
  NOR2XL U336 ( .A(n385), .B(n383), .Y(n222) );
  NAND2XL U337 ( .A(b_15_), .B(b_2_), .Y(n191) );
  NOR2XL U338 ( .A(n391), .B(n381), .Y(n204) );
  NOR2XL U339 ( .A(n388), .B(n385), .Y(n246) );
  NAND2XL U340 ( .A(b_15_), .B(b_6_), .Y(n187) );
  NOR2XL U341 ( .A(n387), .B(n382), .Y(n212) );
  NOR2XL U342 ( .A(n386), .B(n383), .Y(n223) );
  NOR2XL U343 ( .A(n401), .B(n382), .Y(n214) );
  NAND2XL U344 ( .A(b_15_), .B(b_4_), .Y(n189) );
  NOR2XL U345 ( .A(n388), .B(n383), .Y(n225) );
  NOR2XL U346 ( .A(n387), .B(n383), .Y(n224) );
  NAND2XL U347 ( .A(b_15_), .B(b_5_), .Y(n188) );
  NOR2XL U348 ( .A(n386), .B(n384), .Y(n234) );
  NOR2XL U349 ( .A(n386), .B(n381), .Y(n198) );
  NOR2XL U350 ( .A(n384), .B(n383), .Y(n221) );
  NOR2XL U351 ( .A(n385), .B(n382), .Y(n210) );
  NAND2XL U352 ( .A(b_15_), .B(b_8_), .Y(n185) );
  NAND2XL U353 ( .A(b_15_), .B(b_9_), .Y(n184) );
  NOR2XL U354 ( .A(n385), .B(n381), .Y(n197) );
  NOR2XL U355 ( .A(n384), .B(n382), .Y(n209) );
  NOR2XL U356 ( .A(n382), .B(n381), .Y(n194) );
  NAND2XL U357 ( .A(b_15_), .B(b_12_), .Y(n181) );
  NAND2XL U358 ( .A(b_15_), .B(b_11_), .Y(n182) );
  NOR2XL U359 ( .A(n383), .B(n381), .Y(n195) );
  NOR2XL U360 ( .A(n384), .B(n381), .Y(n196) );
  NAND2XL U361 ( .A(b_15_), .B(b_10_), .Y(n183) );
  NOR2XL U362 ( .A(n383), .B(n382), .Y(n208) );
  ADDFXL U363 ( .A(n32), .B(n31), .CI(n4), .CO(n3), .S(product_28_) );
  ADDFXL U364 ( .A(n38), .B(n36), .CI(n6), .CO(n5), .S(product_26_) );
  INVXL U365 ( .A(b_8_), .Y(n399) );
  INVXL U366 ( .A(b_11_), .Y(n396) );
  INVXL U367 ( .A(b_7_), .Y(n400) );
  INVXL U368 ( .A(b_9_), .Y(n398) );
  INVXL U369 ( .A(b_10_), .Y(n397) );
  INVXL U370 ( .A(b_12_), .Y(n395) );
  INVXL U371 ( .A(b_13_), .Y(n394) );
  INVXL U372 ( .A(b_14_), .Y(n393) );
  CLKBUFX2 U373 ( .A(b_0_), .Y(product_0_) );
  CLKINVX1 U374 ( .A(n1), .Y(product_31_) );
  NOR2X1 U375 ( .A(n392), .B(n405), .Y(n297) );
  NOR2X1 U376 ( .A(n392), .B(n389), .Y(n288) );
  NOR2X1 U377 ( .A(n406), .B(n389), .Y(n287) );
  NOR2X1 U378 ( .A(n392), .B(n401), .Y(n283) );
  NOR2X1 U379 ( .A(n405), .B(n401), .Y(n281) );
  NOR2X1 U380 ( .A(n390), .B(n401), .Y(n279) );
  NOR2X1 U381 ( .A(n389), .B(n401), .Y(n278) );
  NOR2X1 U382 ( .A(n392), .B(n388), .Y(n277) );
  NOR2X1 U383 ( .A(n406), .B(n388), .Y(n276) );
  NOR2X1 U384 ( .A(n405), .B(n388), .Y(n275) );
  NOR2X1 U385 ( .A(n401), .B(n388), .Y(n271) );
  NOR2X1 U386 ( .A(n387), .B(n390), .Y(n266) );
  NOR2X1 U387 ( .A(n387), .B(n389), .Y(n265) );
  NOR2X1 U388 ( .A(n387), .B(n401), .Y(n264) );
  NOR2X1 U389 ( .A(n392), .B(n386), .Y(n262) );
  NOR2X1 U390 ( .A(n406), .B(n386), .Y(n261) );
  NOR2X1 U391 ( .A(n405), .B(n386), .Y(n260) );
  NOR2X1 U392 ( .A(n390), .B(n386), .Y(n258) );
  NOR2X1 U393 ( .A(n389), .B(n386), .Y(n257) );
  NOR2X1 U394 ( .A(n401), .B(n386), .Y(n256) );
  NOR2X1 U395 ( .A(n388), .B(n386), .Y(n255) );
  NOR2X1 U396 ( .A(n387), .B(n386), .Y(n254) );
  NOR2X1 U397 ( .A(n392), .B(n385), .Y(n253) );
  NOR2X1 U398 ( .A(n405), .B(n385), .Y(n251) );
  NOR2X1 U399 ( .A(n390), .B(n385), .Y(n249) );
  NOR2X1 U400 ( .A(n401), .B(n385), .Y(n247) );
  NOR2X1 U401 ( .A(n387), .B(n385), .Y(n245) );
  NOR2X1 U402 ( .A(n392), .B(n384), .Y(n243) );
  NOR2X1 U403 ( .A(n406), .B(n384), .Y(n242) );
  NOR2X1 U404 ( .A(n405), .B(n384), .Y(n241) );
  NOR2X1 U405 ( .A(n390), .B(n384), .Y(n239) );
  NOR2X1 U406 ( .A(n389), .B(n384), .Y(n238) );
  NOR2X1 U407 ( .A(n401), .B(n384), .Y(n237) );
  NOR2X1 U408 ( .A(n388), .B(n384), .Y(n236) );
  NOR2X1 U409 ( .A(n385), .B(n384), .Y(n233) );
  NOR2X1 U410 ( .A(n392), .B(n383), .Y(n232) );
  NOR2X1 U411 ( .A(n405), .B(n383), .Y(n230) );
  NOR2X1 U412 ( .A(n389), .B(n383), .Y(n227) );
  NOR2X1 U413 ( .A(n401), .B(n383), .Y(n226) );
  NOR2X1 U414 ( .A(n392), .B(n382), .Y(n220) );
  NOR2X1 U415 ( .A(n406), .B(n382), .Y(n219) );
  NOR2X1 U416 ( .A(n405), .B(n382), .Y(n218) );
  NOR2X1 U417 ( .A(n390), .B(n382), .Y(n216) );
  NOR2X1 U418 ( .A(n389), .B(n382), .Y(n215) );
  NOR2X1 U419 ( .A(n388), .B(n382), .Y(n213) );
  NOR2X1 U420 ( .A(n386), .B(n382), .Y(n211) );
  NOR2X1 U421 ( .A(n392), .B(n381), .Y(n207) );
  NOR2X1 U422 ( .A(n390), .B(n381), .Y(n203) );
  NOR2X1 U423 ( .A(n389), .B(n381), .Y(n202) );
  NOR2X1 U424 ( .A(n401), .B(n381), .Y(n201) );
  NOR2X1 U425 ( .A(n388), .B(n381), .Y(n200) );
endmodule


module Analysis_shift_1mux_DW01_add_0 ( SUM, A_31_, A_30_, A_29_, A_28_, A_27_, 
        A_26_, A_25_, A_24_, A_23_, A_22_, A_21_, A_20_, A_19_, A_18_, A_17_, 
        A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, 
        A_6_, A_5_, A_4_, A_3_, A_2_, A_0_, B_31_, B_30_, B_29_, B_28_, B_27_, 
        B_26_, B_25_, B_24_, B_23_, B_22_, B_21_, B_20_, B_19_, B_18_, B_17_, 
        B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_0_ );
  output [31:0] SUM;
  input A_31_, A_30_, A_29_, A_28_, A_27_, A_26_, A_25_, A_24_, A_23_, A_22_,
         A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_0_,
         B_31_, B_30_, B_29_, B_28_, B_27_, B_26_, B_25_, B_24_, B_23_, B_22_,
         B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_,
         B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_0_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [31:4] carry;

  ADDFX2 U1_29 ( .A(A_29_), .B(B_29_), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_27 ( .A(A_27_), .B(B_27_), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_25 ( .A(A_25_), .B(B_25_), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_23 ( .A(A_23_), .B(B_23_), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX1 U1_3 ( .A(A_3_), .B(B_3_), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X2 U1_31 ( .A(A_31_), .B(B_31_), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFHX1 U1_26 ( .A(A_26_), .B(B_26_), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX1 U1_24 ( .A(A_24_), .B(B_24_), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFHX1 U1_28 ( .A(A_28_), .B(B_28_), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFHX1 U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFHX1 U1_20 ( .A(A_20_), .B(B_20_), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFHX1 U1_22 ( .A(A_22_), .B(B_22_), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFHX2 U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFHX2 U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFHX2 U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFHX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFHX4 U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFHX4 U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFHX4 U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFHX2 U1_30 ( .A(A_30_), .B(B_30_), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  NAND3X2 U1 ( .A(n5), .B(n6), .C(n7), .Y(carry[9]) );
  NAND3X1 U2 ( .A(n2), .B(n3), .C(n4), .Y(carry[12]) );
  NAND2X1 U3 ( .A(B_11_), .B(carry[11]), .Y(n2) );
  AND2X2 U4 ( .A(B_2_), .B(A_2_), .Y(n1) );
  XOR3XL U5 ( .A(carry[11]), .B(A_11_), .C(B_11_), .Y(SUM[11]) );
  NAND2X2 U6 ( .A(A_11_), .B(carry[11]), .Y(n3) );
  NAND2X1 U7 ( .A(A_11_), .B(B_11_), .Y(n4) );
  NAND2X1 U8 ( .A(B_8_), .B(carry[8]), .Y(n5) );
  NAND2X1 U9 ( .A(A_8_), .B(carry[8]), .Y(n6) );
  XOR3XL U10 ( .A(carry[8]), .B(A_8_), .C(B_8_), .Y(SUM[8]) );
  NAND2X1 U11 ( .A(A_8_), .B(B_8_), .Y(n7) );
  NAND2X1 U12 ( .A(B_15_), .B(carry[15]), .Y(n8) );
  NAND2X1 U13 ( .A(A_15_), .B(carry[15]), .Y(n9) );
  NAND2X1 U14 ( .A(A_15_), .B(B_15_), .Y(n10) );
  NAND3X1 U15 ( .A(n8), .B(n9), .C(n10), .Y(carry[16]) );
  XOR3XL U16 ( .A(carry[15]), .B(A_15_), .C(B_15_), .Y(SUM[15]) );
  XOR2XL U17 ( .A(B_2_), .B(A_2_), .Y(SUM[2]) );
  XOR2X1 U18 ( .A(B_0_), .B(A_0_), .Y(SUM[0]) );
  AND2X2 U19 ( .A(B_0_), .B(A_0_), .Y(SUM[1]) );
endmodule


module Analysis_shift_1mux ( clk, rst, fft_valid, fft_d0, done, freq );
  input [31:0] fft_d0;
  output [3:0] freq;
  input clk, rst, fft_valid;
  output done;
  wire   n112, n113, n114, n115, N10, N11, N12, N13, N18, N25, n6, n8, n1100,
         n120, n130, n14, n17, n180, n19, n20, n21, n22, n23, n24, n250, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         mul_out_9_, mul_out_8_, mul_out_7_, mul_out_6_, mul_out_5_,
         mul_out_4_, mul_out_3_, mul_out_31_, mul_out_30_, mul_out_2_,
         mul_out_29_, mul_out_28_, mul_out_27_, mul_out_26_, mul_out_25_,
         mul_out_24_, mul_out_23_, mul_out_22_, mul_out_21_, mul_out_20_,
         mul_out_19_, mul_out_18_, mul_out_17_, mul_out_16_, mul_out_15_,
         mul_out_14_, mul_out_13_, mul_out_12_, mul_out_11_, mul_out_10_,
         mul_out_0_, mul_out2_9_, mul_out2_8_, mul_out2_7_, mul_out2_6_,
         mul_out2_5_, mul_out2_4_, mul_out2_3_, mul_out2_31_, mul_out2_30_,
         mul_out2_2_, mul_out2_29_, mul_out2_28_, mul_out2_27_, mul_out2_26_,
         mul_out2_25_, mul_out2_24_, mul_out2_23_, mul_out2_22_, mul_out2_21_,
         mul_out2_20_, mul_out2_19_, mul_out2_18_, mul_out2_17_, mul_out2_16_,
         mul_out2_15_, mul_out2_14_, mul_out2_13_, mul_out2_12_, mul_out2_11_,
         mul_out2_10_, mul_out2_0_, n3, n4, n16, n87, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n1101;
  wire   [31:0] all_squr;
  wire   [31:0] mux_in2;
  wire   [3:0] compare_result_num;

  Analysis_shift_1mux_DW_cmp_0 gte_935 ( .A(mux_in2), .B(all_squr), 
        .GE_LT_GT_LE(N18) );
  Analysis_shift_1mux_DW_mult_uns_1 mult_929 ( .a_15_(fft_d0[31]), .a_14_(
        fft_d0[30]), .a_13_(fft_d0[29]), .a_12_(fft_d0[28]), .a_11_(fft_d0[27]), .a_10_(fft_d0[26]), .a_9_(fft_d0[25]), .a_7_(fft_d0[23]), .a_6_(fft_d0[22]), 
        .a_5_(fft_d0[21]), .a_4_(fft_d0[20]), .a_3_(fft_d0[19]), .a_2_(
        fft_d0[18]), .a_1_(fft_d0[17]), .b_15_(fft_d0[31]), .b_14_(fft_d0[30]), 
        .b_13_(fft_d0[29]), .b_12_(fft_d0[28]), .b_11_(fft_d0[27]), .b_10_(
        fft_d0[26]), .b_9_(fft_d0[25]), .b_8_(fft_d0[24]), .b_7_(fft_d0[23]), 
        .b_6_(fft_d0[22]), .b_5_(fft_d0[21]), .b_4_(fft_d0[20]), .b_3_(
        fft_d0[19]), .b_2_(fft_d0[18]), .b_1_(fft_d0[17]), .b_0_(fft_d0[16]), 
        .product_31_(mul_out2_31_), .product_30_(mul_out2_30_), .product_29_(
        mul_out2_29_), .product_28_(mul_out2_28_), .product_27_(mul_out2_27_), 
        .product_26_(mul_out2_26_), .product_25_(mul_out2_25_), .product_24_(
        mul_out2_24_), .product_23_(mul_out2_23_), .product_22_(mul_out2_22_), 
        .product_21_(mul_out2_21_), .product_20_(mul_out2_20_), .product_19_(
        mul_out2_19_), .product_18_(mul_out2_18_), .product_17_(mul_out2_17_), 
        .product_16_(mul_out2_16_), .product_15_(mul_out2_15_), .product_14_(
        mul_out2_14_), .product_13_(mul_out2_13_), .product_12_(mul_out2_12_), 
        .product_11_(mul_out2_11_), .product_10_(mul_out2_10_), .product_9_(
        mul_out2_9_), .product_8_(mul_out2_8_), .product_7_(mul_out2_7_), 
        .product_6_(mul_out2_6_), .product_5_(mul_out2_5_), .product_4_(
        mul_out2_4_), .product_3_(mul_out2_3_), .product_2_(mul_out2_2_), 
        .product_0_(mul_out2_0_) );
  Analysis_shift_1mux_DW_mult_uns_0 mult_927 ( .a_15_(fft_d0[15]), .a_14_(
        fft_d0[14]), .a_13_(fft_d0[13]), .a_12_(fft_d0[12]), .a_11_(fft_d0[11]), .a_10_(fft_d0[10]), .a_9_(fft_d0[9]), .a_7_(fft_d0[7]), .a_6_(fft_d0[6]), 
        .a_5_(fft_d0[5]), .a_4_(fft_d0[4]), .a_3_(fft_d0[3]), .a_2_(fft_d0[2]), 
        .a_1_(fft_d0[1]), .b_15_(fft_d0[15]), .b_14_(fft_d0[14]), .b_13_(
        fft_d0[13]), .b_12_(fft_d0[12]), .b_11_(fft_d0[11]), .b_10_(fft_d0[10]), .b_9_(fft_d0[9]), .b_8_(fft_d0[8]), .b_7_(fft_d0[7]), .b_6_(fft_d0[6]), 
        .b_5_(fft_d0[5]), .b_4_(fft_d0[4]), .b_3_(fft_d0[3]), .b_2_(fft_d0[2]), 
        .b_1_(fft_d0[1]), .b_0_(fft_d0[0]), .product_31_(mul_out_31_), 
        .product_30_(mul_out_30_), .product_29_(mul_out_29_), .product_28_(
        mul_out_28_), .product_27_(mul_out_27_), .product_26_(mul_out_26_), 
        .product_25_(mul_out_25_), .product_24_(mul_out_24_), .product_23_(
        mul_out_23_), .product_22_(mul_out_22_), .product_21_(mul_out_21_), 
        .product_20_(mul_out_20_), .product_19_(mul_out_19_), .product_18_(
        mul_out_18_), .product_17_(mul_out_17_), .product_16_(mul_out_16_), 
        .product_15_(mul_out_15_), .product_14_(mul_out_14_), .product_13_(
        mul_out_13_), .product_12_(mul_out_12_), .product_11_(mul_out_11_), 
        .product_10_(mul_out_10_), .product_9_(mul_out_9_), .product_8_(
        mul_out_8_), .product_7_(mul_out_7_), .product_6_(mul_out_6_), 
        .product_5_(mul_out_5_), .product_4_(mul_out_4_), .product_3_(
        mul_out_3_), .product_2_(mul_out_2_), .product_0_(mul_out_0_) );
  Analysis_shift_1mux_DW01_add_0 add_930 ( .SUM(all_squr), .A_31_(mul_out_31_), 
        .A_30_(mul_out_30_), .A_29_(mul_out_29_), .A_28_(mul_out_28_), .A_27_(
        mul_out_27_), .A_26_(mul_out_26_), .A_25_(mul_out_25_), .A_24_(
        mul_out_24_), .A_23_(mul_out_23_), .A_22_(mul_out_22_), .A_21_(
        mul_out_21_), .A_20_(mul_out_20_), .A_19_(mul_out_19_), .A_18_(
        mul_out_18_), .A_17_(mul_out_17_), .A_16_(mul_out_16_), .A_15_(
        mul_out_15_), .A_14_(mul_out_14_), .A_13_(mul_out_13_), .A_12_(
        mul_out_12_), .A_11_(mul_out_11_), .A_10_(mul_out_10_), .A_9_(
        mul_out_9_), .A_8_(mul_out_8_), .A_7_(mul_out_7_), .A_6_(mul_out_6_), 
        .A_5_(mul_out_5_), .A_4_(mul_out_4_), .A_3_(mul_out_3_), .A_2_(
        mul_out_2_), .A_0_(mul_out_0_), .B_31_(mul_out2_31_), .B_30_(
        mul_out2_30_), .B_29_(mul_out2_29_), .B_28_(mul_out2_28_), .B_27_(
        mul_out2_27_), .B_26_(mul_out2_26_), .B_25_(mul_out2_25_), .B_24_(
        mul_out2_24_), .B_23_(mul_out2_23_), .B_22_(mul_out2_22_), .B_21_(
        mul_out2_21_), .B_20_(mul_out2_20_), .B_19_(mul_out2_19_), .B_18_(
        mul_out2_18_), .B_17_(mul_out2_17_), .B_16_(mul_out2_16_), .B_15_(
        mul_out2_15_), .B_14_(mul_out2_14_), .B_13_(mul_out2_13_), .B_12_(
        mul_out2_12_), .B_11_(mul_out2_11_), .B_10_(mul_out2_10_), .B_9_(
        mul_out2_9_), .B_8_(mul_out2_8_), .B_7_(mul_out2_7_), .B_6_(
        mul_out2_6_), .B_5_(mul_out2_5_), .B_4_(mul_out2_4_), .B_3_(
        mul_out2_3_), .B_2_(mul_out2_2_), .B_0_(mul_out2_0_) );
  DFFRX1 cnt_state_reg ( .D(n96), .CK(clk), .RN(n1101), .QN(n180) );
  DFFRX1 comp_max_reg_0_ ( .D(n86), .CK(clk), .RN(n1101), .Q(mux_in2[0]), .QN(
        n54) );
  DFFRX1 comp_max_reg_31_ ( .D(n85), .CK(clk), .RN(n98), .Q(mux_in2[31]), .QN(
        n53) );
  DFFRX1 comp_max_reg_30_ ( .D(n84), .CK(clk), .RN(n98), .Q(mux_in2[30]), .QN(
        n52) );
  DFFRX1 comp_max_reg_26_ ( .D(n80), .CK(clk), .RN(n98), .Q(mux_in2[26]), .QN(
        n48) );
  DFFRX1 comp_max_reg_24_ ( .D(n78), .CK(clk), .RN(n98), .Q(mux_in2[24]), .QN(
        n46) );
  DFFRX1 comp_max_reg_20_ ( .D(n74), .CK(clk), .RN(n98), .Q(mux_in2[20]), .QN(
        n42) );
  DFFRX1 comp_max_reg_18_ ( .D(n72), .CK(clk), .RN(n97), .Q(mux_in2[18]), .QN(
        n40) );
  DFFRX1 comp_max_reg_6_ ( .D(n60), .CK(clk), .RN(n87), .Q(mux_in2[6]), .QN(
        n28) );
  DFFRX1 comp_max_reg_4_ ( .D(n58), .CK(clk), .RN(n87), .Q(mux_in2[4]), .QN(
        n26) );
  DFFRX1 comp_max_reg_1_ ( .D(n55), .CK(clk), .RN(n87), .Q(mux_in2[1]), .QN(
        n23) );
  DFFRX1 comp_max_reg_28_ ( .D(n82), .CK(clk), .RN(n98), .Q(mux_in2[28]), .QN(
        n50) );
  DFFRX1 comp_max_reg_16_ ( .D(n70), .CK(clk), .RN(n97), .Q(mux_in2[16]), .QN(
        n38) );
  DFFRX1 comp_max_reg_27_ ( .D(n81), .CK(clk), .RN(n98), .Q(mux_in2[27]), .QN(
        n49) );
  DFFRX1 comp_max_reg_25_ ( .D(n79), .CK(clk), .RN(n98), .Q(mux_in2[25]), .QN(
        n47) );
  DFFRX1 comp_max_reg_23_ ( .D(n77), .CK(clk), .RN(n98), .Q(mux_in2[23]), .QN(
        n45) );
  DFFRX1 comp_max_reg_22_ ( .D(n76), .CK(clk), .RN(n98), .Q(mux_in2[22]), .QN(
        n44) );
  DFFRX1 comp_max_reg_21_ ( .D(n75), .CK(clk), .RN(n98), .Q(mux_in2[21]), .QN(
        n43) );
  DFFRX1 comp_max_reg_19_ ( .D(n73), .CK(clk), .RN(n97), .Q(mux_in2[19]), .QN(
        n41) );
  DFFRX1 comp_max_reg_15_ ( .D(n69), .CK(clk), .RN(n97), .Q(mux_in2[15]), .QN(
        n37) );
  DFFRX1 comp_max_reg_14_ ( .D(n68), .CK(clk), .RN(n97), .Q(mux_in2[14]), .QN(
        n36) );
  DFFRX1 comp_max_reg_7_ ( .D(n61), .CK(clk), .RN(n87), .Q(mux_in2[7]), .QN(
        n29) );
  DFFRX1 comp_max_reg_29_ ( .D(n83), .CK(clk), .RN(n98), .Q(mux_in2[29]), .QN(
        n51) );
  DFFRX1 comp_max_reg_17_ ( .D(n71), .CK(clk), .RN(n97), .Q(mux_in2[17]), .QN(
        n39) );
  DFFRX1 comp_max_reg_13_ ( .D(n67), .CK(clk), .RN(n97), .Q(mux_in2[13]), .QN(
        n35) );
  DFFRX1 comp_max_reg_11_ ( .D(n65), .CK(clk), .RN(n97), .Q(mux_in2[11]), .QN(
        n33) );
  DFFRX1 comp_max_reg_9_ ( .D(n63), .CK(clk), .RN(n97), .Q(mux_in2[9]), .QN(
        n31) );
  DFFRX1 comp_max_reg_3_ ( .D(n57), .CK(clk), .RN(n87), .Q(mux_in2[3]), .QN(
        n250) );
  DFFRX1 comp_max_reg_10_ ( .D(n64), .CK(clk), .RN(n97), .Q(mux_in2[10]), .QN(
        n32) );
  DFFRX1 comp_max_reg_2_ ( .D(n56), .CK(clk), .RN(n87), .Q(mux_in2[2]), .QN(
        n24) );
  DFFRX1 comp_max_reg_12_ ( .D(n66), .CK(clk), .RN(n97), .Q(mux_in2[12]), .QN(
        n34) );
  DFFRX1 comp_max_reg_8_ ( .D(n62), .CK(clk), .RN(n97), .Q(mux_in2[8]), .QN(
        n30) );
  DFFRX1 comp_max_reg_5_ ( .D(n59), .CK(clk), .RN(n87), .Q(mux_in2[5]), .QN(
        n27) );
  DFFRX1 cnt_reg_1_ ( .D(N11), .CK(clk), .RN(n97), .QN(n90) );
  DFFRX1 cnt_reg_0_ ( .D(N10), .CK(clk), .RN(n87), .QN(n91) );
  DFFRX1 cnt_reg_2_ ( .D(N12), .CK(clk), .RN(n98), .Q(n3), .QN(n89) );
  DFFRX1 cnt_reg_3_ ( .D(N13), .CK(clk), .RN(n87), .QN(n88) );
  DFFQX1 freq_reg_0_ ( .D(compare_result_num[0]), .CK(clk), .Q(n115) );
  DFFRX2 compare_result_num_reg_0_ ( .D(n92), .CK(clk), .RN(n87), .Q(
        compare_result_num[0]), .QN(n22) );
  DFFQX1 freq_reg_1_ ( .D(compare_result_num[1]), .CK(clk), .Q(n114) );
  DFFRX2 compare_result_num_reg_1_ ( .D(n93), .CK(clk), .RN(n87), .Q(
        compare_result_num[1]), .QN(n21) );
  DFFQX1 freq_reg_2_ ( .D(compare_result_num[2]), .CK(clk), .Q(n113) );
  DFFRX2 compare_result_num_reg_2_ ( .D(n94), .CK(clk), .RN(n87), .Q(
        compare_result_num[2]), .QN(n20) );
  DFFQX1 freq_reg_3_ ( .D(compare_result_num[3]), .CK(clk), .Q(n112) );
  DFFRHQX1 done_reg ( .D(N25), .CK(clk), .RN(n1101), .Q(n16) );
  DFFRX1 compare_result_num_reg_3_ ( .D(n95), .CK(clk), .RN(n87), .Q(
        compare_result_num[3]), .QN(n19) );
  INVX12 U3 ( .A(n105), .Y(n99) );
  INVX20 U4 ( .A(n103), .Y(n102) );
  INVX8 U7 ( .A(n104), .Y(n101) );
  OAI2BB2X2 U8 ( .B0(n34), .B1(n100), .A0N(all_squr[12]), .A1N(n101), .Y(n66)
         );
  INVX6 U9 ( .A(n104), .Y(n100) );
  CLKBUFX3 U10 ( .A(n106), .Y(n104) );
  OAI2BB2XL U11 ( .B0(n24), .B1(n101), .A0N(all_squr[2]), .A1N(n102), .Y(n56)
         );
  OAI2BB2XL U12 ( .B0(n250), .B1(n101), .A0N(all_squr[3]), .A1N(n102), .Y(n57)
         );
  OAI2BB2XL U13 ( .B0(n31), .B1(n101), .A0N(all_squr[9]), .A1N(n102), .Y(n63)
         );
  OAI2BB2XL U14 ( .B0(n23), .B1(n101), .A0N(all_squr[1]), .A1N(n102), .Y(n55)
         );
  OAI2BB2XL U15 ( .B0(n26), .B1(n101), .A0N(all_squr[4]), .A1N(n102), .Y(n58)
         );
  INVXL U16 ( .A(n16), .Y(n4) );
  INVX12 U17 ( .A(n4), .Y(done) );
  BUFX3 U18 ( .A(n106), .Y(n103) );
  BUFX12 U19 ( .A(n112), .Y(freq[3]) );
  BUFX12 U20 ( .A(n113), .Y(freq[2]) );
  BUFX12 U21 ( .A(n114), .Y(freq[1]) );
  BUFX12 U22 ( .A(n115), .Y(freq[0]) );
  OAI22XL U23 ( .A0(n19), .A1(n101), .B0(n88), .B1(n106), .Y(n95) );
  INVX4 U24 ( .A(n6), .Y(n106) );
  NAND2X2 U25 ( .A(N18), .B(n8), .Y(n6) );
  CLKINVX1 U26 ( .A(rst), .Y(n1101) );
  CLKBUFX3 U27 ( .A(n106), .Y(n105) );
  CLKINVX1 U28 ( .A(n14), .Y(n107) );
  NAND2X1 U29 ( .A(n14), .B(n108), .Y(n17) );
  CLKINVX1 U30 ( .A(n130), .Y(n108) );
  CLKBUFX3 U31 ( .A(n1101), .Y(n87) );
  CLKBUFX3 U32 ( .A(n1101), .Y(n97) );
  CLKBUFX3 U33 ( .A(n1101), .Y(n98) );
  OAI22XL U34 ( .A0(n89), .A1(n105), .B0(n20), .B1(n101), .Y(n94) );
  OAI22XL U35 ( .A0(n90), .A1(n105), .B0(n21), .B1(n101), .Y(n93) );
  OAI22XL U36 ( .A0(n91), .A1(n105), .B0(n22), .B1(n101), .Y(n92) );
  OAI2BB2XL U37 ( .B0(n27), .B1(n100), .A0N(all_squr[5]), .A1N(n102), .Y(n59)
         );
  OAI2BB2XL U38 ( .B0(n28), .B1(n101), .A0N(all_squr[6]), .A1N(n102), .Y(n60)
         );
  OAI2BB2XL U39 ( .B0(n29), .B1(n101), .A0N(all_squr[7]), .A1N(n102), .Y(n61)
         );
  OAI2BB2XL U40 ( .B0(n30), .B1(n101), .A0N(all_squr[8]), .A1N(n102), .Y(n62)
         );
  OAI2BB2XL U41 ( .B0(n32), .B1(n100), .A0N(all_squr[10]), .A1N(n102), .Y(n64)
         );
  OAI2BB2XL U42 ( .B0(n33), .B1(n100), .A0N(all_squr[11]), .A1N(n102), .Y(n65)
         );
  OAI2BB2XL U43 ( .B0(n35), .B1(n100), .A0N(all_squr[13]), .A1N(n102), .Y(n67)
         );
  OAI2BB2XL U44 ( .B0(n36), .B1(n100), .A0N(all_squr[14]), .A1N(n102), .Y(n68)
         );
  OAI2BB2XL U45 ( .B0(n37), .B1(n100), .A0N(all_squr[15]), .A1N(n102), .Y(n69)
         );
  OAI2BB2XL U46 ( .B0(n38), .B1(n100), .A0N(all_squr[16]), .A1N(n102), .Y(n70)
         );
  OAI2BB2XL U47 ( .B0(n39), .B1(n100), .A0N(all_squr[17]), .A1N(n102), .Y(n71)
         );
  OAI2BB2XL U48 ( .B0(n40), .B1(n100), .A0N(all_squr[18]), .A1N(n102), .Y(n72)
         );
  OAI2BB2XL U49 ( .B0(n41), .B1(n100), .A0N(all_squr[19]), .A1N(n102), .Y(n73)
         );
  OAI2BB2XL U50 ( .B0(n42), .B1(n100), .A0N(all_squr[20]), .A1N(n102), .Y(n74)
         );
  OAI2BB2XL U51 ( .B0(n43), .B1(n99), .A0N(all_squr[21]), .A1N(n102), .Y(n75)
         );
  OAI2BB2XL U52 ( .B0(n44), .B1(n99), .A0N(all_squr[22]), .A1N(n102), .Y(n76)
         );
  OAI2BB2XL U53 ( .B0(n45), .B1(n99), .A0N(all_squr[23]), .A1N(n102), .Y(n77)
         );
  OAI2BB2XL U54 ( .B0(n46), .B1(n99), .A0N(all_squr[24]), .A1N(n102), .Y(n78)
         );
  OAI2BB2XL U55 ( .B0(n47), .B1(n99), .A0N(all_squr[25]), .A1N(n102), .Y(n79)
         );
  OAI2BB2XL U56 ( .B0(n48), .B1(n99), .A0N(all_squr[26]), .A1N(n102), .Y(n80)
         );
  OAI2BB2XL U57 ( .B0(n49), .B1(n99), .A0N(all_squr[27]), .A1N(n102), .Y(n81)
         );
  OAI2BB2XL U58 ( .B0(n50), .B1(n99), .A0N(all_squr[28]), .A1N(n102), .Y(n82)
         );
  OAI2BB2XL U59 ( .B0(n51), .B1(n99), .A0N(all_squr[29]), .A1N(n102), .Y(n83)
         );
  OAI2BB2XL U60 ( .B0(n52), .B1(n99), .A0N(all_squr[30]), .A1N(n102), .Y(n84)
         );
  OAI2BB2XL U61 ( .B0(n53), .B1(n99), .A0N(all_squr[31]), .A1N(n102), .Y(n85)
         );
  OAI2BB2XL U62 ( .B0(n54), .B1(n99), .A0N(all_squr[0]), .A1N(n102), .Y(n86)
         );
  NAND4X1 U63 ( .A(n88), .B(n89), .C(n90), .D(n91), .Y(n8) );
  INVXL U64 ( .A(fft_valid), .Y(n109) );
  OAI32X1 U65 ( .A0(n108), .A1(n107), .A2(n3), .B0(n89), .B1(n17), .Y(N12) );
  NAND2X1 U66 ( .A(n180), .B(n109), .Y(n14) );
  AOI211X1 U67 ( .A0(n90), .A1(n91), .B0(n107), .C0(n130), .Y(N11) );
  OAI21XL U68 ( .A0(n1100), .A1(n88), .B0(n120), .Y(N13) );
  NAND4X1 U69 ( .A(n130), .B(n88), .C(n14), .D(n3), .Y(n120) );
  OA21XL U70 ( .A0(n107), .A1(n3), .B0(n17), .Y(n1100) );
  NOR2BX1 U71 ( .AN(n91), .B(n107), .Y(N10) );
  OAI21XL U72 ( .A0(n180), .A1(N25), .B0(n109), .Y(n96) );
  NOR3X1 U73 ( .A(n89), .B(n88), .C(n108), .Y(N25) );
  NOR2X1 U74 ( .A(n91), .B(n90), .Y(n130) );
endmodule


module FAS ( data_valid, data, clk, rst, fir_d, fir_valid, fft_valid, done, 
        freq, fft_d1, fft_d2, fft_d3, fft_d4, fft_d5, fft_d6, fft_d7, fft_d8, 
        fft_d9, fft_d10, fft_d11, fft_d12, fft_d13, fft_d14, fft_d15, fft_d0
 );
  input [15:0] data;
  output [15:0] fir_d;
  output [3:0] freq;
  output [31:0] fft_d1;
  output [31:0] fft_d2;
  output [31:0] fft_d3;
  output [31:0] fft_d4;
  output [31:0] fft_d5;
  output [31:0] fft_d6;
  output [31:0] fft_d7;
  output [31:0] fft_d8;
  output [31:0] fft_d9;
  output [31:0] fft_d10;
  output [31:0] fft_d11;
  output [31:0] fft_d12;
  output [31:0] fft_d13;
  output [31:0] fft_d14;
  output [31:0] fft_d15;
  output [31:0] fft_d0;
  input data_valid, clk, rst;
  output fir_valid, fft_valid, done;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n2, n4, n6, n8, n10, n12, n14, n16, n18, n20, n22, n24, n26,
         n28, n30;

  FIR_FILTER2 fir_filter0 ( .clk(clk), .rst(rst), .data_valid(data_valid), 
        .data(data), .fir_valid(fir_valid), .fir_d(fir_d) );
  FFT_ultrafast2_shift FFT0 ( .clk(clk), .rst(rst), .fir_valid(fir_valid), 
        .fir_d(fir_d), .fft_valid(fft_valid), .fft_d1(fft_d1), .fft_d2(fft_d2), 
        .fft_d3(fft_d3), .fft_d4(fft_d4), .fft_d5(fft_d5), .fft_d6(fft_d6), 
        .fft_d7(fft_d7), .fft_d8(fft_d8), .fft_d9(fft_d9), .fft_d10(fft_d10), 
        .fft_d11(fft_d11), .fft_d12(fft_d12), .fft_d13(fft_d13), .fft_d14(
        fft_d14), .fft_d15(fft_d15), .fft_d0({fft_d0[31:26], n32, n33, n34, 
        fft_d0[22], n35, n36, fft_d0[19], n37, n38, fft_d0[16:12], n39, 
        fft_d0[10], n40, n41, n42, fft_d0[6], n43, n44, n45, n46, n47, 
        fft_d0[0]}) );
  Analysis_shift_1mux Analysis0 ( .clk(clk), .rst(rst), .fft_valid(fft_valid), 
        .fft_d0(fft_d0), .done(done), .freq(freq) );
  CLKBUFX20 U1 ( .A(n39), .Y(fft_d0[11]) );
  INVX12 U2 ( .A(n32), .Y(n2) );
  CLKINVX20 U3 ( .A(n2), .Y(fft_d0[25]) );
  INVX12 U4 ( .A(n40), .Y(n4) );
  CLKINVX20 U5 ( .A(n4), .Y(fft_d0[9]) );
  INVX12 U6 ( .A(n34), .Y(n6) );
  CLKINVX20 U7 ( .A(n6), .Y(fft_d0[23]) );
  INVX12 U8 ( .A(n33), .Y(n8) );
  CLKINVX20 U9 ( .A(n8), .Y(fft_d0[24]) );
  INVX12 U10 ( .A(n41), .Y(n10) );
  CLKINVX20 U11 ( .A(n10), .Y(fft_d0[8]) );
  CLKINVX20 U12 ( .A(n26), .Y(fft_d0[21]) );
  INVX8 U13 ( .A(n42), .Y(n12) );
  CLKINVX20 U14 ( .A(n12), .Y(fft_d0[7]) );
  CLKINVX20 U15 ( .A(n18), .Y(fft_d0[2]) );
  CLKINVX20 U16 ( .A(n16), .Y(fft_d0[18]) );
  INVX8 U17 ( .A(n45), .Y(n14) );
  CLKINVX20 U18 ( .A(n14), .Y(fft_d0[3]) );
  INVX3 U19 ( .A(n46), .Y(n18) );
  INVX3 U20 ( .A(n37), .Y(n16) );
  INVX3 U21 ( .A(n35), .Y(n26) );
  CLKINVX12 U22 ( .A(n47), .Y(n20) );
  CLKINVX20 U23 ( .A(n20), .Y(fft_d0[1]) );
  CLKINVX12 U24 ( .A(n38), .Y(n22) );
  CLKINVX20 U25 ( .A(n22), .Y(fft_d0[17]) );
  CLKINVX12 U26 ( .A(n43), .Y(n24) );
  CLKINVX20 U27 ( .A(n24), .Y(fft_d0[5]) );
  CLKINVX12 U28 ( .A(n44), .Y(n28) );
  CLKINVX20 U29 ( .A(n28), .Y(fft_d0[4]) );
  CLKINVX12 U30 ( .A(n36), .Y(n30) );
  CLKINVX20 U31 ( .A(n30), .Y(fft_d0[20]) );
endmodule

